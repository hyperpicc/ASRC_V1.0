library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package src_rom_pkg is

	constant COE_WIDTH	: integer := 26;
	constant COE_CENTRE	: signed( 25 downto 0 ) := b"01111111010111000010100100";

	type COE_ROM_TYPE is array( 4095 downto 0 ) of signed( 25 downto 0 );
	constant COE_ROM	 : COE_ROM_TYPE := (
		b"01111111010110010001101101",
		b"01111111010011111111001000",
		b"01111111010000001010111001",
		b"01111111001010110101000110",
		b"01111111000011111101110101",
		b"01111110111011100101010000",
		b"01111110110001101011100011",
		b"01111110100110010000111011",
		b"01111110011001010101101000",
		b"01111110001010111001111100",
		b"01111101111010111110001100",
		b"01111101101001100010101100",
		b"01111101010110100111110110",
		b"01111101000010001110000011",
		b"01111100101100010101110000",
		b"01111100010100111111011011",
		b"01111011111100001011100011",
		b"01111011100001111010101101",
		b"01111011000110001101011011",
		b"01111010101001000100010011",
		b"01111010001010100000000000",
		b"01111001101010100001001001",
		b"01111001001001001000011100",
		b"01111000100110010110100110",
		b"01111000000010001100011000",
		b"01110111011100101010100011",
		b"01110110110101110001111010",
		b"01110110001101100011010100",
		b"01110101100011111111100111",
		b"01110100111001000111101101",
		b"01110100001100111100100000",
		b"01110011011111011110111101",
		b"01110010110000110000000010",
		b"01110010000000110000110000",
		b"01110001001111100010000111",
		b"01110000011101000101001100",
		b"01101111101001011011000011",
		b"01101110110100100100110011",
		b"01101101111110100011100011",
		b"01101101000111011000011110",
		b"01101100001111000100101110",
		b"01101011010101101001011111",
		b"01101010011011001000000001",
		b"01101001011111100001100011",
		b"01101000100010110111010100",
		b"01100111100101001010101000",
		b"01100110100110011100110010",
		b"01100101100110101111000111",
		b"01100100100110000010111011",
		b"01100011100100011001101000",
		b"01100010100001110100100101",
		b"01100001011110010101001011",
		b"01100000011001111100110101",
		b"01011111010100101100111111",
		b"01011110001110100111000110",
		b"01011101000111101100101000",
		b"01011011111111111111000010",
		b"01011010110111011111110101",
		b"01011001101110010000100001",
		b"01011000100100010010100111",
		b"01010111011001100111101010",
		b"01010110001110010001001101",
		b"01010101000010010000110010",
		b"01010011110101100111111111",
		b"01010010101000011000011001",
		b"01010001011010100011100100",
		b"01010000001100001011001000",
		b"01001110111101010000101010",
		b"01001101101101110101110011",
		b"01001100011101111100001001",
		b"01001011001101100101010101",
		b"01001001111100110011000000",
		b"01001000101011100110110001",
		b"01000111011010000010010010",
		b"01000110001000000111001101",
		b"01000100110101110111001010",
		b"01000011100011010011110100",
		b"01000010010000011110110100",
		b"01000000111101011001110100",
		b"00111111101010000110011110",
		b"00111110010110100110011101",
		b"00111101000010111011011001",
		b"00111011101111000110111101",
		b"00111010011011001010110010",
		b"00111001000111001000100010",
		b"00110111110011000001110111",
		b"00110110011110111000011001",
		b"00110101001010101101110001",
		b"00110011110110100011101000",
		b"00110010100010011011100110",
		b"00110001001110010111010010",
		b"00101111111010011000010101",
		b"00101110100110100000010100",
		b"00101101010010110000110110",
		b"00101011111111001011100001",
		b"00101010101011110001111011",
		b"00101001011000100101100110",
		b"00101000000101101000001001",
		b"00100110110010111011000101",
		b"00100101100000011111111101",
		b"00100100001110011000010011",
		b"00100010111100100101100111",
		b"00100001101011001001011010",
		b"00100000011010000101001100",
		b"00011111001001011010011001",
		b"00011101111001001010011111",
		b"00011100101001010110111011",
		b"00011011011010000001001000",
		b"00011010001011001010100000",
		b"00011000111100110100011100",
		b"00010111101111000000010100",
		b"00010110100001101111100000",
		b"00010101010101000011010100",
		b"00010100001000111101000101",
		b"00010010111101011110000111",
		b"00010001110010100111101100",
		b"00010000101000011011000100",
		b"00001111011110111001011110",
		b"00001110010110000100001010",
		b"00001101001101111100010010",
		b"00001100000110100011000011",
		b"00001010111111111001100111",
		b"00001001111010000001000101",
		b"00001000110100111010100101",
		b"00000111110000100111001100",
		b"00000110101101000111111111",
		b"00000101101010011101111110",
		b"00000100101000101010001100",
		b"00000011100111101101100111",
		b"00000010100111101001001110",
		b"00000001101000011101111011",
		b"00000000101010001100101010",
		b"11111111101100110110010011",
		b"11111110110000011011101101",
		b"11111101110100111101101101",
		b"11111100111010011101001000",
		b"11111100000000111010101111",
		b"11111011001000010111010001",
		b"11111010010000110011011110",
		b"11111001011010010000000011",
		b"11111000100100101101101010",
		b"11110111110000001100111100",
		b"11110110111100101110100000",
		b"11110110001010010010111101",
		b"11110101011000111010110110",
		b"11110100101000100110101100",
		b"11110011111001010111000000",
		b"11110011001011001100010001",
		b"11110010011110000110111010",
		b"11110001110010000111010110",
		b"11110001000111001101111110",
		b"11110000011101011011001000",
		b"11101111110100101111001011",
		b"11101111001101001010011000",
		b"11101110100110101101000010",
		b"11101110000001010111011000",
		b"11101101011101001001101000",
		b"11101100111010000011111100",
		b"11101100011000000110100000",
		b"11101011110111010001011100",
		b"11101011010111100100110101",
		b"11101010111001000000110001",
		b"11101010011011100101010010",
		b"11101001111111010010011000",
		b"11101001100100001000000011",
		b"11101001001010000110010000",
		b"11101000110001001100111011",
		b"11101000011001011011111100",
		b"11101000000010110011001101",
		b"11100111101101010010100010",
		b"11100111011000111001110001",
		b"11100111000101101000101100",
		b"11100110110011011111000100",
		b"11100110100010011100101000",
		b"11100110010010100001000101",
		b"11100110000011101100001000",
		b"11100101110101111101011011",
		b"11100101101001010100100101",
		b"11100101011101110001001110",
		b"11100101010011010010111011",
		b"11100101001001111001010000",
		b"11100101000001100011101111",
		b"11100100111010010001111000",
		b"11100100110100000011001010",
		b"11100100101110110111000011",
		b"11100100101010101100111111",
		b"11100100100111100100011000",
		b"11100100100101011100100111",
		b"11100100100100010101000011",
		b"11100100100100001101000100",
		b"11100100100101000011111110",
		b"11100100100110111001000100",
		b"11100100101001101011101000",
		b"11100100101101011010111100",
		b"11100100110010000110001110",
		b"11100100110111101100101110",
		b"11100100111110001101101000",
		b"11100101000101101000001000",
		b"11100101001101111011011001",
		b"11100101010111000110100100",
		b"11100101100001001000110010",
		b"11100101101100000001001010",
		b"11100101110111101110110011",
		b"11100110000100010000110010",
		b"11100110010001100110001011",
		b"11100110011111101110000010",
		b"11100110101110100111011001",
		b"11100110111110010001010001",
		b"11100111001110101010101100",
		b"11100111011111110010101000",
		b"11100111110001101000000110",
		b"11101000000100001010000011",
		b"11101000010111010111011100",
		b"11101000101011001111001111",
		b"11101000111111110000011000",
		b"11101001010100111001110010",
		b"11101001101010101010011000",
		b"11101010000001000001000100",
		b"11101010010111111100110000",
		b"11101010101111011100010110",
		b"11101011000111011110101101",
		b"11101011100000000010101111",
		b"11101011111001000111010011",
		b"11101100010010101011010001",
		b"11101100101100101101100000",
		b"11101101000111001100110111",
		b"11101101100010001000001100",
		b"11101101111101011110010110",
		b"11101110011001001110001010",
		b"11101110110101010110100000",
		b"11101111010001110110001100",
		b"11101111101110101100000101",
		b"11110000001011110111000000",
		b"11110000101001010101110011",
		b"11110001000111000111010100",
		b"11110001100101001010010111",
		b"11110010000011011101110011",
		b"11110010100010000000011110",
		b"11110011000000110001001101",
		b"11110011011111101110110110",
		b"11110011111110111000010001",
		b"11110100011110001100010011",
		b"11110100111101101001110011",
		b"11110101011101001111101000",
		b"11110101111100111100101001",
		b"11110110011100101111101110",
		b"11110110111100100111110000",
		b"11110111011100100011100111",
		b"11110111111100100010001010",
		b"11111000011100100010010101",
		b"11111000111100100011000001",
		b"11111001011100100011001000",
		b"11111001111100100001100101",
		b"11111010011100011101010100",
		b"11111010111100010101010001",
		b"11111011011100001000011000",
		b"11111011111011110101101000",
		b"11111100011011011011111110",
		b"11111100111010111010011001",
		b"11111101011010001111111000",
		b"11111101111001011011011101",
		b"11111110011000011100001000",
		b"11111110110111010000111100",
		b"11111111010101111000111010",
		b"11111111110100010011001000",
		b"00000000010010011110101000",
		b"00000000110000011010100010",
		b"00000001001110000101111010",
		b"00000001101011011111111010",
		b"00000010001000100111101000",
		b"00000010100101011100001111",
		b"00000011000001111100111000",
		b"00000011011110001000110000",
		b"00000011111001111111000010",
		b"00000100010101011110111100",
		b"00000100110000100111101100",
		b"00000101001011011000100011",
		b"00000101100101110000110001",
		b"00000101111111101111101000",
		b"00000110011001010100011100",
		b"00000110110010011110100000",
		b"00000111001011001101001001",
		b"00000111100011011111110000",
		b"00000111111011010101101010",
		b"00001000010010101110010010",
		b"00001000101001101001000010",
		b"00001001000000000101010101",
		b"00001001010110000010101001",
		b"00001001101011100000011010",
		b"00001010000000011110001000",
		b"00001010010100111011010101",
		b"00001010101000110111100001",
		b"00001010111100010010010001",
		b"00001011001111001011000111",
		b"00001011100001100001101011",
		b"00001011110011010101100011",
		b"00001100000100100110010111",
		b"00001100010101010011110001",
		b"00001100100101011101011101",
		b"00001100110101000011000110",
		b"00001101000100000100011010",
		b"00001101010010100001000111",
		b"00001101100000011001000000",
		b"00001101101101101011110100",
		b"00001101111010011001010110",
		b"00001110000110100001011100",
		b"00001110010010000011111010",
		b"00001110011101000000100111",
		b"00001110100111010111011100",
		b"00001110110001001000010010",
		b"00001110111010010011000100",
		b"00001111000010110111101101",
		b"00001111001010110110001100",
		b"00001111010010001110011110",
		b"00001111011001000000100100",
		b"00001111011111001100011111",
		b"00001111100100110010010010",
		b"00001111101001110001111111",
		b"00001111101110001011101101",
		b"00001111110001111111100001",
		b"00001111110101001101100011",
		b"00001111110111110101111011",
		b"00001111111001111000110011",
		b"00001111111011010110010111",
		b"00001111111100001110110001",
		b"00001111111100100010010001",
		b"00001111111100010001000100",
		b"00001111111011011011011010",
		b"00001111111010000001100100",
		b"00001111111000000011110011",
		b"00001111110101100010011100",
		b"00001111110010011101110001",
		b"00001111101110110110000111",
		b"00001111101010101011110110",
		b"00001111100101111111010100",
		b"00001111100000110000111010",
		b"00001111011011000001000000",
		b"00001111010100110000000001",
		b"00001111001101111110011000",
		b"00001111000110101100100001",
		b"00001110111110111010111001",
		b"00001110110110101001111110",
		b"00001110101101111010001111",
		b"00001110100100101100001010",
		b"00001110011011000000010010",
		b"00001110010000110111000111",
		b"00001110000110010001001010",
		b"00001101111011001111000000",
		b"00001101101111110001001010",
		b"00001101100011111000001111",
		b"00001101010111100100110010",
		b"00001101001010110111011010",
		b"00001100111101110000101100",
		b"00001100110000010001010000",
		b"00001100100010011001101101",
		b"00001100010100001010101011",
		b"00001100000101100100110100",
		b"00001011110110101000110000",
		b"00001011100111010111001001",
		b"00001011010111110000101010",
		b"00001011000111110101111101",
		b"00001010110111100111101101",
		b"00001010100111000110100110",
		b"00001010010110010011010100",
		b"00001010000101001110100011",
		b"00001001110011111001000000",
		b"00001001100010010011011000",
		b"00001001010000011110011001",
		b"00001000111110011010101111",
		b"00001000101100001001001001",
		b"00001000011001101010010101",
		b"00001000000110111111000000",
		b"00000111110100000111111010",
		b"00000111100001000101110001",
		b"00000111001101111001010011",
		b"00000110111010100011001111",
		b"00000110100111000100010101",
		b"00000110010011011101010010",
		b"00000101111111101110110111",
		b"00000101101011111001110000",
		b"00000101010111111110101111",
		b"00000101000011111110100000",
		b"00000100101111111001110100",
		b"00000100011011110001011000",
		b"00000100000111100101111100",
		b"00000011110011011000001100",
		b"00000011011111001000111001",
		b"00000011001010111000101110",
		b"00000010110110101000011011",
		b"00000010100010011000101101",
		b"00000010001110001010010001",
		b"00000001111001111101110100",
		b"00000001100101110100000010",
		b"00000001010001101101101000",
		b"00000000111101101011010010",
		b"00000000101001101101101100",
		b"00000000010101110101100000",
		b"00000000000010000011011010",
		b"11111111101110011000000011",
		b"11111111011010110100000110",
		b"11111111000111011000001100",
		b"11111110110100000100111110",
		b"11111110100000111011000100",
		b"11111110001101111011000111",
		b"11111101111011000101101101",
		b"11111101101000011011011110",
		b"11111101010101111100111111",
		b"11111101000011101010110110",
		b"11111100110001100101101000",
		b"11111100011111101101111001",
		b"11111100001110000100001110",
		b"11111011111100101001001000",
		b"11111011101011011101001011",
		b"11111011011010100000110111",
		b"11111011001001110100101110",
		b"11111010111001011001010001",
		b"11111010101001001110111110",
		b"11111010011001010110010011",
		b"11111010001001101111110000",
		b"11111001111010011011110001",
		b"11111001101011011010110011",
		b"11111001011100101101010000",
		b"11111001001110010011100101",
		b"11111001000000001110001010",
		b"11111000110010011101011001",
		b"11111000100101000001101011",
		b"11111000010111111011010101",
		b"11111000001011001010110000",
		b"11110111111110110000010001",
		b"11110111110010101100001100",
		b"11110111100110111110110110",
		b"11110111011011101000100010",
		b"11110111010000101001100001",
		b"11110111000110000010000101",
		b"11110110111011110010011111",
		b"11110110110001111010111110",
		b"11110110101000011011110000",
		b"11110110011111010101000011",
		b"11110110010110100111000100",
		b"11110110001110010001111111",
		b"11110110000110010101111110",
		b"11110101111110110011001100",
		b"11110101110111101001110001",
		b"11110101110000111001110110",
		b"11110101101010100011100010",
		b"11110101100100100110111011",
		b"11110101011111000100000110",
		b"11110101011001111011001001",
		b"11110101010101001100000110",
		b"11110101010000110111000000",
		b"11110101001100111011111001",
		b"11110101001001011010110001",
		b"11110101000110010011101001",
		b"11110101000011100110100000",
		b"11110101000001010011010011",
		b"11110100111111011001111111",
		b"11110100111101111010100010",
		b"11110100111100110100110110",
		b"11110100111100001000110110",
		b"11110100111011110110011011",
		b"11110100111011111101100000",
		b"11110100111100011101111010",
		b"11110100111101010111100010",
		b"11110100111110101010001110",
		b"11110101000000010101110100",
		b"11110101000010011010000111",
		b"11110101000100110110111100",
		b"11110101000111101100000110",
		b"11110101001010111001011000",
		b"11110101001110011110100010",
		b"11110101010010011011010101",
		b"11110101010110101111100010",
		b"11110101011011011010110111",
		b"11110101100000011101000011",
		b"11110101100101110101110100",
		b"11110101101011100100110111",
		b"11110101110001101001111001",
		b"11110101111000000100100100",
		b"11110101111110110100100101",
		b"11110110000101111001100101",
		b"11110110001101010011001111",
		b"11110110010101000001001011",
		b"11110110011101000011000010",
		b"11110110100101011000011100",
		b"11110110101110000001000000",
		b"11110110110110111100010110",
		b"11110111000000001010000011",
		b"11110111001001101001101101",
		b"11110111010011011010111011",
		b"11110111011101011101001111",
		b"11110111100111110000001111",
		b"11110111110010010011011111",
		b"11110111111101000110100001",
		b"11111000001000001000111010",
		b"11111000010011011010001010",
		b"11111000011110111001110110",
		b"11111000101010100111011110",
		b"11111000110110100010100011",
		b"11111001000010101010101000",
		b"11111001001110111111001101",
		b"11111001011011011111110010",
		b"11111001101000001011110111",
		b"11111001110101000010111101",
		b"11111010000010000100100011",
		b"11111010001111010000001001",
		b"11111010011100100101001110",
		b"11111010101010000011010001",
		b"11111010110111101001110010",
		b"11111011000101011000001110",
		b"11111011010011001110000100",
		b"11111011100001001010110100",
		b"11111011101111001101111011",
		b"11111011111101010110110111",
		b"11111100001011100101001000",
		b"11111100011001111000001100",
		b"11111100101000001111100000",
		b"11111100110110101010100010",
		b"11111101000101001000110010",
		b"11111101010011101001101101",
		b"11111101100010001100110010",
		b"11111101110000110001100000",
		b"11111101111111010111010011",
		b"11111110001101111101101100",
		b"11111110011100100100001001",
		b"11111110101011001010001001",
		b"11111110111001101111001011",
		b"11111111001000010010101101",
		b"11111111010110110100010000",
		b"11111111100101010011010011",
		b"11111111110011101111010110",
		b"00000000000010000111111001",
		b"00000000010000011100011100",
		b"00000000011110101100011111",
		b"00000000101100110111100100",
		b"00000000111010111101001100",
		b"00000001001000111100111001",
		b"00000001010110110110001011",
		b"00000001100100101000100110",
		b"00000001110010010011101100",
		b"00000001111111110111000000",
		b"00000010001101010010000100",
		b"00000010011010100100011110",
		b"00000010100111101101110001",
		b"00000010110100101101100010",
		b"00000011000001100011010101",
		b"00000011001110001110110000",
		b"00000011011010101111011010",
		b"00000011100111000100111001",
		b"00000011110011001110110011",
		b"00000011111111001100110000",
		b"00000100001010111110011000",
		b"00000100010110100011010100",
		b"00000100100001111011001101",
		b"00000100101101000101101100",
		b"00000100111000000010011100",
		b"00000101000010110001000110",
		b"00000101001101010001011000",
		b"00000101010111100010111100",
		b"00000101100001100101011111",
		b"00000101101011011000101110",
		b"00000101110100111100010111",
		b"00000101111110010000001001",
		b"00000110000111010011110010",
		b"00000110010000000111000010",
		b"00000110011000101001101001",
		b"00000110100000111011011000",
		b"00000110101000111100000001",
		b"00000110110000101011010110",
		b"00000110111000001001001010",
		b"00000110111111010101010000",
		b"00000111000110001111011101",
		b"00000111001100110111100110",
		b"00000111010011001101100000",
		b"00000111011001010001000001",
		b"00000111011111000010000001",
		b"00000111100100100000010111",
		b"00000111101001101011111100",
		b"00000111101110100100101000",
		b"00000111110011001010010110",
		b"00000111110111011100111111",
		b"00000111111011011100011111",
		b"00000111111111001000110001",
		b"00001000000010100001110011",
		b"00001000000101100111100001",
		b"00001000001000011001111001",
		b"00001000001010111000111010",
		b"00001000001101000100100011",
		b"00001000001110111100110101",
		b"00001000010000100001101110",
		b"00001000010001110011010010",
		b"00001000010010110001100010",
		b"00001000010011011100100000",
		b"00001000010011110100010001",
		b"00001000010011111000110111",
		b"00001000010011101010011000",
		b"00001000010011001000111000",
		b"00001000010010010100011111",
		b"00001000010001001101010010",
		b"00001000001111110011011001",
		b"00001000001110000110111011",
		b"00001000001100001000000001",
		b"00001000001001110110110101",
		b"00001000000111010011011111",
		b"00001000000100011110001011",
		b"00001000000001010111000010",
		b"00000111111101111110010010",
		b"00000111111010010100000101",
		b"00000111110110011000101000",
		b"00000111110010001100001001",
		b"00000111101101101110110101",
		b"00000111101001000000111011",
		b"00000111100100000010101010",
		b"00000111011110110100010000",
		b"00000111011001010101111110",
		b"00000111010011101000000011",
		b"00000111001101101010110010",
		b"00000111000111011110011011",
		b"00000111000001000011010000",
		b"00000110111010011001100011",
		b"00000110110011100001100111",
		b"00000110101100011011101111",
		b"00000110100101001000001111",
		b"00000110011101100111011010",
		b"00000110010101111001100101",
		b"00000110001101111111000101",
		b"00000110000101111000001110",
		b"00000101111101100101010111",
		b"00000101110101000110110100",
		b"00000101101100011100111101",
		b"00000101100011101000000111",
		b"00000101011010101000101010",
		b"00000101010001011110111100",
		b"00000101001000001011010100",
		b"00000100111110101110001011",
		b"00000100110101000111111000",
		b"00000100101011011000110011",
		b"00000100100001100001010100",
		b"00000100010111100001110100",
		b"00000100001101011010101100",
		b"00000100000011001100010100",
		b"00000011111000110111000110",
		b"00000011101110011011011010",
		b"00000011100011111001101010",
		b"00000011011001010010001111",
		b"00000011001110100101100100",
		b"00000011000011110100000000",
		b"00000010111000111101111111",
		b"00000010101110000011111010",
		b"00000010100011000110001011",
		b"00000010011000000101001011",
		b"00000010001101000001010101",
		b"00000010000001111011000010",
		b"00000001110110110010101101",
		b"00000001101011101000101110",
		b"00000001100000011101100001",
		b"00000001010101010001011110",
		b"00000001001010000100111111",
		b"00000000111110111000011110",
		b"00000000110011101100010101",
		b"00000000101000100000111100",
		b"00000000011101010110101110",
		b"00000000010010001110000011",
		b"00000000000111000111010101",
		b"11111111111100000010111011",
		b"11111111110001000001010000",
		b"11111111100110000010101010",
		b"11111111011011000111100100",
		b"11111111010000010000010100",
		b"11111111000101011101010011",
		b"11111110111010101110111000",
		b"11111110110000000101011011",
		b"11111110100101100001010011",
		b"11111110011011000010110110",
		b"11111110010000101010011011",
		b"11111110000110011000011001",
		b"11111101111100001101000110",
		b"11111101110010001000110110",
		b"11111101101000001100000000",
		b"11111101011110010110111000",
		b"11111101010100101001110011",
		b"11111101001011000101000110",
		b"11111101000001101001000011",
		b"11111100111000010110000000",
		b"11111100101111001100001110",
		b"11111100100110001100000001",
		b"11111100011101010101101011",
		b"11111100010100101001011101",
		b"11111100001100000111101010",
		b"11111100000011110000100011",
		b"11111011111011100100011000",
		b"11111011110011100011011001",
		b"11111011101011101101110110",
		b"11111011100100000011111110",
		b"11111011011100100110000000",
		b"11111011010101010100001011",
		b"11111011001110001110101100",
		b"11111011000111010101110001",
		b"11111011000000101001100110",
		b"11111010111010001010011000",
		b"11111010110011111000010011",
		b"11111010101101110011100010",
		b"11111010100111111100010001",
		b"11111010100010010010101000",
		b"11111010011100110110110010",
		b"11111010010111101000111001",
		b"11111010010010101001000110",
		b"11111010001101110111011111",
		b"11111010001001010100001110",
		b"11111010000100111111011001",
		b"11111010000000111001000111",
		b"11111001111101000001011110",
		b"11111001111001011000100100",
		b"11111001110101111110011110",
		b"11111001110010110011001111",
		b"11111001101111110110111101",
		b"11111001101101001001101010",
		b"11111001101010101011011001",
		b"11111001101000011100001101",
		b"11111001100110011100000111",
		b"11111001100100101011001001",
		b"11111001100011001001010011",
		b"11111001100001110110100101",
		b"11111001100000110010111111",
		b"11111001011111111110100000",
		b"11111001011111011001000111",
		b"11111001011111000010110001",
		b"11111001011110111011011101",
		b"11111001011111000011000110",
		b"11111001011111011001101010",
		b"11111001011111111111000100",
		b"11111001100000110011010000",
		b"11111001100001110110001001",
		b"11111001100011000111101000",
		b"11111001100100100111101000",
		b"11111001100110010110000011",
		b"11111001101000010010110001",
		b"11111001101010011101101011",
		b"11111001101100110110101000",
		b"11111001101111011101100000",
		b"11111001110010010010001010",
		b"11111001110101010100011101",
		b"11111001111000100100001111",
		b"11111001111100000001010101",
		b"11111001111111101011100100",
		b"11111010000011100010110010",
		b"11111010000111100110110011",
		b"11111010001011110111011010",
		b"11111010010000010100011100",
		b"11111010010100111101101011",
		b"11111010011001110010111010",
		b"11111010011110110011111100",
		b"11111010100100000000100010",
		b"11111010101001011000011110",
		b"11111010101110111011100010",
		b"11111010110100101001011110",
		b"11111010111010100010000011",
		b"11111011000000100101000010",
		b"11111011000110110010001001",
		b"11111011001101001001001010",
		b"11111011010011101001110010",
		b"11111011011010010011110010",
		b"11111011100001000110111001",
		b"11111011101000000010110011",
		b"11111011101111000111010001",
		b"11111011110110010100000000",
		b"11111011111101101000101101",
		b"11111100000101000101000111",
		b"11111100001100101000111010",
		b"11111100010100010011110100",
		b"11111100011100000101100010",
		b"11111100100011111101110001",
		b"11111100101011111100001101",
		b"11111100110100000000100010",
		b"11111100111100001010011110",
		b"11111101000100011001101100",
		b"11111101001100101101111000",
		b"11111101010101000110101110",
		b"11111101011101100011111011",
		b"11111101100110000101001001",
		b"11111101101110101010000101",
		b"11111101110111010010011010",
		b"11111101111111111101110100",
		b"11111110001000101011111110",
		b"11111110010001011100100100",
		b"11111110011010001111010001",
		b"11111110100011000011110010",
		b"11111110101011111001110000",
		b"11111110110100110000111000",
		b"11111110111101101000110110",
		b"11111111000110100001010100",
		b"11111111001111011001111111",
		b"11111111011000010010100010",
		b"11111111100001001010101001",
		b"11111111101010000010000000",
		b"11111111110010111000010010",
		b"11111111111011101101001100",
		b"00000000000100100000011001",
		b"00000000001101010001100111",
		b"00000000010110000000100001",
		b"00000000011110101100110100",
		b"00000000100111010110001101",
		b"00000000101111111100011001",
		b"00000000111000011111000011",
		b"00000001000000111101111011",
		b"00000001001001011000101101",
		b"00000001010001101111000111",
		b"00000001011010000000110110",
		b"00000001100010001101101001",
		b"00000001101010010101001111",
		b"00000001110010010111010100",
		b"00000001111010010011101010",
		b"00000010000010001001111101",
		b"00000010001001111001111111",
		b"00000010010001100011011110",
		b"00000010011001000110001010",
		b"00000010100000100001110011",
		b"00000010100111110110001011",
		b"00000010101111000011000001",
		b"00000010110110001000000111",
		b"00000010111101000101001110",
		b"00000011000011111010001001",
		b"00000011001010100110101000",
		b"00000011010001001010011111",
		b"00000011010111100101100000",
		b"00000011011101110111011111",
		b"00000011100100000000001111",
		b"00000011101001111111100100",
		b"00000011101111110101010010",
		b"00000011110101100001001110",
		b"00000011111011000011001100",
		b"00000100000000011011000011",
		b"00000100000101101000101000",
		b"00000100001010101011110001",
		b"00000100001111100100010101",
		b"00000100010100010010001010",
		b"00000100011000110101001001",
		b"00000100011101001101001001",
		b"00000100100001011010000011",
		b"00000100100101011011101110",
		b"00000100101001010010000101",
		b"00000100101100111101000000",
		b"00000100110000011100011010",
		b"00000100110011110000001100",
		b"00000100110110111000010011",
		b"00000100111001110100101000",
		b"00000100111100100101001000",
		b"00000100111111001001101111",
		b"00000101000001100010011001",
		b"00000101000011101111000011",
		b"00000101000101101111101011",
		b"00000101000111100100001110",
		b"00000101001001001100101100",
		b"00000101001010101001000001",
		b"00000101001011111001001111",
		b"00000101001100111101010100",
		b"00000101001101110101010000",
		b"00000101001110100001000100",
		b"00000101001111000000110000",
		b"00000101001111010100010111",
		b"00000101001111011011111001",
		b"00000101001111010111011001",
		b"00000101001111000110111001",
		b"00000101001110101010011101",
		b"00000101001110000010001000",
		b"00000101001101001101111101",
		b"00000101001100001110000010",
		b"00000101001011000010011001",
		b"00000101001001101011001010",
		b"00000101001000001000011001",
		b"00000101000110011010001011",
		b"00000101000100100000101000",
		b"00000101000010011011110110",
		b"00000101000000001011111011",
		b"00000100111101110000111111",
		b"00000100111011001011001010",
		b"00000100111000011010100100",
		b"00000100110101011111010110",
		b"00000100110010011001101000",
		b"00000100101111001001100011",
		b"00000100101011101111010001",
		b"00000100101000001010111011",
		b"00000100100100011100101101",
		b"00000100100000100100110000",
		b"00000100011100100011001110",
		b"00000100011000011000010100",
		b"00000100010100000100001101",
		b"00000100001111100111000100",
		b"00000100001011000001000101",
		b"00000100000110010010011101",
		b"00000100000001011011011000",
		b"00000011111100011100000010",
		b"00000011110111010100101010",
		b"00000011110010000101011011",
		b"00000011101100101110100101",
		b"00000011100111010000010011",
		b"00000011100001101010110101",
		b"00000011011011111110011001",
		b"00000011010110001011001100",
		b"00000011010000010001011110",
		b"00000011001010010001011110",
		b"00000011000100001011011001",
		b"00000010111101111111100000",
		b"00000010110111101110000010",
		b"00000010110001010111001110",
		b"00000010101010111011010011",
		b"00000010100100011010100010",
		b"00000010011101110101001010",
		b"00000010010111001011011100",
		b"00000010010000011101100110",
		b"00000010001001101011111010",
		b"00000010000010110110101000",
		b"00000001111011111101111111",
		b"00000001110101000010010001",
		b"00000001101110000011101110",
		b"00000001100111000010100110",
		b"00000001011111111111001001",
		b"00000001011000111001101001",
		b"00000001010001110010010110",
		b"00000001001010101001100001",
		b"00000001000011011111011010",
		b"00000000111100010100010010",
		b"00000000110101001000011001",
		b"00000000101101111100000000",
		b"00000000100110101111010111",
		b"00000000011111100010110000",
		b"00000000011000010110011010",
		b"00000000010001001010100110",
		b"00000000001001111111100100",
		b"00000000000010110101100100",
		b"11111111111011101100110111",
		b"11111111110100100101101101",
		b"11111111101101100000010101",
		b"11111111100110011100111111",
		b"11111111011111011011111011",
		b"11111111011000011101011001",
		b"11111111010001100001101001",
		b"11111111001010101000111000",
		b"11111111000011110011011000",
		b"11111110111101000001010101",
		b"11111110110110010011000001",
		b"11111110101111101000101000",
		b"11111110101001000010011010",
		b"11111110100010100000100100",
		b"11111110011100000011010110",
		b"11111110010101101010111100",
		b"11111110001111010111100100",
		b"11111110001001001001011100",
		b"11111110000011000000110001",
		b"11111101111100111101110000",
		b"11111101110111000000100110",
		b"11111101110001001001011111",
		b"11111101101011011000100111",
		b"11111101100101101110001011",
		b"11111101100000001010010101",
		b"11111101011010101101010011",
		b"11111101010101010111001101",
		b"11111101010000001000010000",
		b"11111101001011000000100111",
		b"11111101000110000000011010",
		b"11111101000001000111110101",
		b"11111100111100010111000001",
		b"11111100110111101110001000",
		b"11111100110011001101010010",
		b"11111100101110110100101000",
		b"11111100101010100100010011",
		b"11111100100110011100011011",
		b"11111100100010011101000111",
		b"11111100011110100110100000",
		b"11111100011010111000101100",
		b"11111100010111010011110010",
		b"11111100010011110111111000",
		b"11111100010000100101000110",
		b"11111100001101011011011111",
		b"11111100001010011011001011",
		b"11111100000111100100001101",
		b"11111100000100110110101011",
		b"11111100000010010010101010",
		b"11111011111111111000001100",
		b"11111011111101100111010110",
		b"11111011111011100000001100",
		b"11111011111001100010101111",
		b"11111011110111101111000100",
		b"11111011110110000101001011",
		b"11111011110100100101000111",
		b"11111011110011001110111010",
		b"11111011110010000010100100",
		b"11111011110001000000000111",
		b"11111011110000000111100011",
		b"11111011101111011000111000",
		b"11111011101110110100000111",
		b"11111011101110011001001101",
		b"11111011101110001000001011",
		b"11111011101110000000111111",
		b"11111011101110000011101000",
		b"11111011101110010000000011",
		b"11111011101110100110001111",
		b"11111011101111000110001000",
		b"11111011101111101111101100",
		b"11111011110000100010110111",
		b"11111011110001011111100110",
		b"11111011110010100101110101",
		b"11111011110011110101011111",
		b"11111011110101001110100000",
		b"11111011110110110000110011",
		b"11111011111000011100010010",
		b"11111011111010010000111000",
		b"11111011111100001110100000",
		b"11111011111110010101000010",
		b"11111100000000100100011001",
		b"11111100000010111100011101",
		b"11111100000101011101001000",
		b"11111100001000000110010010",
		b"11111100001010110111110100",
		b"11111100001101110001100101",
		b"11111100010000110011011110",
		b"11111100010011111101010110",
		b"11111100010111001111000100",
		b"11111100011010101000011111",
		b"11111100011110001001011110",
		b"11111100100001110001111000",
		b"11111100100101100001100011",
		b"11111100101001011000010101",
		b"11111100101101010110000100",
		b"11111100110001011010100101",
		b"11111100110101100101101110",
		b"11111100111001110111010101",
		b"11111100111110001111001101",
		b"11111101000010101101001101",
		b"11111101000111010001001000",
		b"11111101001011111010110011",
		b"11111101010000101010000010",
		b"11111101010101011110101010",
		b"11111101011010011000011110",
		b"11111101011111010111010011",
		b"11111101100100011010111100",
		b"11111101101001100011001100",
		b"11111101101110101111110111",
		b"11111101110100000000110000",
		b"11111101111001010101101011",
		b"11111101111110101110011010",
		b"11111110000100001010110000",
		b"11111110001001101010100001",
		b"11111110001111001101011111",
		b"11111110010100110011011101",
		b"11111110011010011100001101",
		b"11111110100000000111100011",
		b"11111110100101110101010000",
		b"11111110101011100101000111",
		b"11111110110001010110111011",
		b"11111110110111001010011110",
		b"11111110111100111111100011",
		b"11111111000010110101111011",
		b"11111111001000101101011010",
		b"11111111001110100101110001",
		b"11111111010100011110110011",
		b"11111111011010011000010011",
		b"11111111100000010010000010",
		b"11111111100110001011110100",
		b"11111111101100000101011011",
		b"11111111110001111110101001",
		b"11111111110111110111010010",
		b"11111111111101101111000111",
		b"00000000000011100101111011",
		b"00000000001001011011100010",
		b"00000000001111001111101110",
		b"00000000010101000010010001",
		b"00000000011010110011000000",
		b"00000000100000100001101110",
		b"00000000100110001110001101",
		b"00000000101011111000010001",
		b"00000000110001011111101101",
		b"00000000110111000100010110",
		b"00000000111100100101111111",
		b"00000001000010000100011100",
		b"00000001000111011111100000",
		b"00000001001100110111000001",
		b"00000001010010001010110011",
		b"00000001010111011010101010",
		b"00000001011100100110011011",
		b"00000001100001101101111010",
		b"00000001100110110000111110",
		b"00000001101011101111011011",
		b"00000001110000101001000110",
		b"00000001110101011101110111",
		b"00000001111010001101100001",
		b"00000001111110110111111100",
		b"00000010000011011100111101",
		b"00000010000111111100011100",
		b"00000010001100010110001111",
		b"00000010010000101010001101",
		b"00000010010100111000001101",
		b"00000010011001000000000111",
		b"00000010011101000001110010",
		b"00000010100000111101000111",
		b"00000010100100110001111110",
		b"00000010101000100000001110",
		b"00000010101100000111110001",
		b"00000010101111101000100000",
		b"00000010110011000010010100",
		b"00000010110110010101000110",
		b"00000010111001100000110001",
		b"00000010111100100101001110",
		b"00000010111111100010010111",
		b"00000011000010011000001000",
		b"00000011000101000110011011",
		b"00000011000111101101001011",
		b"00000011001010001100010011",
		b"00000011001100100011110000",
		b"00000011001110110011011110",
		b"00000011010000111011011000",
		b"00000011010010111011011011",
		b"00000011010100110011100101",
		b"00000011010110100011110010",
		b"00000011011000001100000000",
		b"00000011011001101100001100",
		b"00000011011011000100010101",
		b"00000011011100010100011001",
		b"00000011011101011100010110",
		b"00000011011110011100001100",
		b"00000011011111010011111001",
		b"00000011100000000011011110",
		b"00000011100000101010111010",
		b"00000011100001001010001100",
		b"00000011100001100001010111",
		b"00000011100001110000011001",
		b"00000011100001110111010100",
		b"00000011100001110110001010",
		b"00000011100001101100111100",
		b"00000011100001011011101011",
		b"00000011100001000010011010",
		b"00000011100000100001001011",
		b"00000011011111111000000000",
		b"00000011011111000110111110",
		b"00000011011110001110000110",
		b"00000011011101001101011101",
		b"00000011011100000101000110",
		b"00000011011010110101000100",
		b"00000011011001011101011110",
		b"00000011010111111110010110",
		b"00000011010110010111110001",
		b"00000011010100101001110101",
		b"00000011010010110100101000",
		b"00000011010000111000001101",
		b"00000011001110110100101100",
		b"00000011001100101010001010",
		b"00000011001010011000101101",
		b"00000011001000000000011100",
		b"00000011000101100001011110",
		b"00000011000010111011111001",
		b"00000011000000001111110101",
		b"00000010111101011101011001",
		b"00000010111010100100101100",
		b"00000010110111100101110110",
		b"00000010110100100000111111",
		b"00000010110001010110010000",
		b"00000010101110000101110000",
		b"00000010101010101111101000",
		b"00000010100111010100000000",
		b"00000010100011110011000011",
		b"00000010100000001100110111",
		b"00000010011100100001101000",
		b"00000010011000110001011101",
		b"00000010010100111100100001",
		b"00000010010001000010111101",
		b"00000010001101000100111011",
		b"00000010001001000010100100",
		b"00000010000100111100000100",
		b"00000010000000110001100011",
		b"00000001111100100011001100",
		b"00000001111000010001001010",
		b"00000001110011111011100110",
		b"00000001101111100010101100",
		b"00000001101011000110100110",
		b"00000001100110100111011111",
		b"00000001100010000101100001",
		b"00000001011101100000111000",
		b"00000001011000111001101110",
		b"00000001010100010000001111",
		b"00000001001111100100100101",
		b"00000001001010110110111011",
		b"00000001000110000111011101",
		b"00000001000001010110010110",
		b"00000000111100100011110001",
		b"00000000110111101111111001",
		b"00000000110010111010111001",
		b"00000000101110000100111101",
		b"00000000101001001110001111",
		b"00000000100100010110111100",
		b"00000000011111011111001110",
		b"00000000011010100111010001",
		b"00000000010101101111001111",
		b"00000000010000110111010100",
		b"00000000001011111111101011",
		b"00000000000111001000011111",
		b"00000000000010010001111011",
		b"11111111111101011100001010",
		b"11111111111000100111010110",
		b"11111111110011110011101100",
		b"11111111101111000001010101",
		b"11111111101010010000011100",
		b"11111111100101100001001011",
		b"11111111100000110011101111",
		b"11111111011100001000001111",
		b"11111111010111011110111000",
		b"11111111010010110111110100",
		b"11111111001110010011001011",
		b"11111111001001110001001001",
		b"11111111000101010001111000",
		b"11111111000000110101100000",
		b"11111110111100011100001100",
		b"11111110111000000110000101",
		b"11111110110011110011010100",
		b"11111110101111100100000100",
		b"11111110101011011000011011",
		b"11111110100111010000100101",
		b"11111110100011001100101001",
		b"11111110011111001100101111",
		b"11111110011011010001000001",
		b"11111110010111011001100111",
		b"11111110010011100110101000",
		b"11111110001111111000001100",
		b"11111110001100001110011011",
		b"11111110001000101001011101",
		b"11111110000101001001011001",
		b"11111110000001101110010110",
		b"11111101111110011000011011",
		b"11111101111011000111101110",
		b"11111101110111111100010111",
		b"11111101110100110110011011",
		b"11111101110001110110000000",
		b"11111101101110111011001101",
		b"11111101101100000110000110",
		b"11111101101001010110110010",
		b"11111101100110101101010110",
		b"11111101100100001001110110",
		b"11111101100001101100011000",
		b"11111101011111010100111111",
		b"11111101011101000011110001",
		b"11111101011010111000110001",
		b"11111101011000110100000011",
		b"11111101010110110101101010",
		b"11111101010100111101101011",
		b"11111101010011001100001000",
		b"11111101010001100001000100",
		b"11111101001111111100100001",
		b"11111101001110011110100011",
		b"11111101001101000111001011",
		b"11111101001011110110011011",
		b"11111101001010101100010101",
		b"11111101001001101000111010",
		b"11111101001000101100001100",
		b"11111101000111110110001100",
		b"11111101000111000110111001",
		b"11111101000110011110010101",
		b"11111101000101111100100000",
		b"11111101000101100001011010",
		b"11111101000101001101000011",
		b"11111101000100111111011010",
		b"11111101000100111000011110",
		b"11111101000100111000001110",
		b"11111101000100111110101010",
		b"11111101000101001011110000",
		b"11111101000101011111011110",
		b"11111101000101111001110010",
		b"11111101000110011010101010",
		b"11111101000111000010000100",
		b"11111101000111101111111110",
		b"11111101001000100100010011",
		b"11111101001001011111000010",
		b"11111101001010100000000111",
		b"11111101001011100111011111",
		b"11111101001100110101000110",
		b"11111101001110001000111000",
		b"11111101001111100010110000",
		b"11111101010001000010101100",
		b"11111101010010101000100101",
		b"11111101010100010100011000",
		b"11111101010110000110000000",
		b"11111101010111111101010111",
		b"11111101011001111010011000",
		b"11111101011011111100111110",
		b"11111101011110000101000011",
		b"11111101100000010010100001",
		b"11111101100010100101010011",
		b"11111101100100111101010001",
		b"11111101100111011010010110",
		b"11111101101001111100011011",
		b"11111101101100100011011001",
		b"11111101101111001111001010",
		b"11111101110001111111100111",
		b"11111101110100110100101000",
		b"11111101110111101110000110",
		b"11111101111010101011111010",
		b"11111101111101101101111100",
		b"11111110000000110100000101",
		b"11111110000011111110001100",
		b"11111110000111001100001011",
		b"11111110001010011101111000",
		b"11111110001101110011001100",
		b"11111110010001001011111110",
		b"11111110010100101000000110",
		b"11111110011000000111011100",
		b"11111110011011101001110111",
		b"11111110011111001111001110",
		b"11111110100010110111011001",
		b"11111110100110100010001111",
		b"11111110101010001111100111",
		b"11111110101101111111011000",
		b"11111110110001110001011010",
		b"11111110110101100101100010",
		b"11111110111001011011101001",
		b"11111110111101010011100101",
		b"11111111000001001101001100",
		b"11111111000101001000010110",
		b"11111111001001000100111001",
		b"11111111001101000010101100",
		b"11111111010001000001100111",
		b"11111111010101000001011110",
		b"11111111011001000010001010",
		b"11111111011101000011100001",
		b"11111111100001000101011010",
		b"11111111100101000111101011",
		b"11111111101001001010001011",
		b"11111111101101001100110001",
		b"11111111110001001111010011",
		b"11111111110101010001101001",
		b"11111111111001010011101001",
		b"11111111111101010101001010",
		b"00000000000001010110000011",
		b"00000000000101010110001100",
		b"00000000001001010101011010",
		b"00000000001101010011100101",
		b"00000000010001010000100100",
		b"00000000010101001100001111",
		b"00000000011001000110011100",
		b"00000000011100111111000100",
		b"00000000100000110101111100",
		b"00000000100100101010111110",
		b"00000000101000011110000000",
		b"00000000101100001110111011",
		b"00000000101111111101100101",
		b"00000000110011101001110111",
		b"00000000110111010011101001",
		b"00000000111010111010110100",
		b"00000000111110011111001110",
		b"00000001000010000000110001",
		b"00000001000101011111010110",
		b"00000001001000111010110100",
		b"00000001001100010011000100",
		b"00000001001111101000000000",
		b"00000001010010111001100000",
		b"00000001010110000111011101",
		b"00000001011001010001110001",
		b"00000001011100011000010110",
		b"00000001011111011011000100",
		b"00000001100010011001110110",
		b"00000001100101010100100101",
		b"00000001101000001011001100",
		b"00000001101010111101100101",
		b"00000001101101101011101010",
		b"00000001110000010101010110",
		b"00000001110010111010100011",
		b"00000001110101011011001100",
		b"00000001110111110111001110",
		b"00000001111010001110100001",
		b"00000001111100100001000100",
		b"00000001111110101110110000",
		b"00000010000000110111100001",
		b"00000010000010111011010101",
		b"00000010000100111010000110",
		b"00000010000110110011110010",
		b"00000010001000101000010100",
		b"00000010001010010111101011",
		b"00000010001100000001110001",
		b"00000010001101100110100110",
		b"00000010001111000110000110",
		b"00000010010000100000001110",
		b"00000010010001110100111101",
		b"00000010010011000100010000",
		b"00000010010100001110000110",
		b"00000010010101010010011101",
		b"00000010010110010001010011",
		b"00000010010111001010101000",
		b"00000010010111111110011001",
		b"00000010011000101100100111",
		b"00000010011001010101010001",
		b"00000010011001111000010101",
		b"00000010011010010101110101",
		b"00000010011010101101110000",
		b"00000010011011000000000101",
		b"00000010011011001100110110",
		b"00000010011011010100000011",
		b"00000010011011010101101101",
		b"00000010011011010001110101",
		b"00000010011011001000011011",
		b"00000010011010111001100001",
		b"00000010011010100101001001",
		b"00000010011010001011010100",
		b"00000010011001101100000100",
		b"00000010011001000111011100",
		b"00000010011000011101011110",
		b"00000010010111101110001011",
		b"00000010010110111001100111",
		b"00000010010101111111110101",
		b"00000010010101000000110111",
		b"00000010010011111100110000",
		b"00000010010010110011100101",
		b"00000010010001100101011000",
		b"00000010010000010010001110",
		b"00000010001110111010001001",
		b"00000010001101011101001111",
		b"00000010001011111011100011",
		b"00000010001010010101001010",
		b"00000010001000101010000111",
		b"00000010000110111010100001",
		b"00000010000101000110011011",
		b"00000010000011001101111010",
		b"00000010000001010001000100",
		b"00000001111111001111111110",
		b"00000001111101001010101101",
		b"00000001111011000001010111",
		b"00000001111000110100000001",
		b"00000001110110100010110001",
		b"00000001110100001101101100",
		b"00000001110001110100111010",
		b"00000001101111011000100000",
		b"00000001101100111000100100",
		b"00000001101010010101001100",
		b"00000001100111101110100000",
		b"00000001100101000100100101",
		b"00000001100010010111100010",
		b"00000001011111100111011110",
		b"00000001011100110100100000",
		b"00000001011001111110101110",
		b"00000001010111000110010000",
		b"00000001010100001011001101",
		b"00000001010001001101101011",
		b"00000001001110001101110010",
		b"00000001001011001011101001",
		b"00000001001000000111011000",
		b"00000001000101000001000110",
		b"00000001000001111000111001",
		b"00000000111110101110111011",
		b"00000000111011100011010010",
		b"00000000111000010110000110",
		b"00000000110101000111011110",
		b"00000000110001110111100010",
		b"00000000101110100110011010",
		b"00000000101011010100001101",
		b"00000000101000000001000011",
		b"00000000100100101101000100",
		b"00000000100001011000010111",
		b"00000000011110000011000100",
		b"00000000011010101101010011",
		b"00000000010111010111001100",
		b"00000000010100000000110101",
		b"00000000010000101010010111",
		b"00000000001101010011111010",
		b"00000000001001111101100101",
		b"00000000000110100111100000",
		b"00000000000011010001110010",
		b"11111111111111111100100010",
		b"11111111111100100111111001",
		b"11111111111001010011111110",
		b"11111111110110000000111000",
		b"11111111110010101110101111",
		b"11111111101111011101101001",
		b"11111111101100001101101111",
		b"11111111101000111111000110",
		b"11111111100101110001111000",
		b"11111111100010100110001001",
		b"11111111011111011100000010",
		b"11111111011100010011101010",
		b"11111111011001001101000111",
		b"11111111010110001000011111",
		b"11111111010011000101111010",
		b"11111111010000000101011110",
		b"11111111001101000111010010",
		b"11111111001010001011011100",
		b"11111111000111010010000010",
		b"11111111000100011011001010",
		b"11111111000001100110111011",
		b"11111110111110110101011010",
		b"11111110111100000110101101",
		b"11111110111001011010111010",
		b"11111110110110110010000111",
		b"11111110110100001100011000",
		b"11111110110001101001110100",
		b"11111110101111001010011111",
		b"11111110101100101110011111",
		b"11111110101010010101111000",
		b"11111110101000000000110000",
		b"11111110100101101111001010",
		b"11111110100011100001001100",
		b"11111110100001010110111011",
		b"11111110011111010000011001",
		b"11111110011101001101101100",
		b"11111110011011001110110110",
		b"11111110011001010011111101",
		b"11111110010111011101000100",
		b"11111110010101101010001110",
		b"11111110010011111011011111",
		b"11111110010010010000111001",
		b"11111110010000101010100001",
		b"11111110001111001000011000",
		b"11111110001101101010100001",
		b"11111110001100010000111111",
		b"11111110001010111011110101",
		b"11111110001001101011000101",
		b"11111110001000011110110000",
		b"11111110000111010110111001",
		b"11111110000110010011100010",
		b"11111110000101010100101011",
		b"11111110000100011010010111",
		b"11111110000011100100100110",
		b"11111110000010110011011010",
		b"11111110000010000110110100",
		b"11111110000001011110110100",
		b"11111110000000111011011100",
		b"11111110000000011100101010",
		b"11111110000000000010100001",
		b"11111101111111101100111111",
		b"11111101111111011100000101",
		b"11111101111111001111110011",
		b"11111101111111001000000111",
		b"11111101111111000101000010",
		b"11111101111111000110100011",
		b"11111101111111001100101001",
		b"11111101111111010111010011",
		b"11111101111111100110011111",
		b"11111101111111111010001101",
		b"11111110000000010010011011",
		b"11111110000000101111000110",
		b"11111110000001010000001110",
		b"11111110000001110101110001",
		b"11111110000010011111101011",
		b"11111110000011001101111100",
		b"11111110000100000000100000",
		b"11111110000100110111010100",
		b"11111110000101110010010111",
		b"11111110000110110001100110",
		b"11111110000111110100111100",
		b"11111110001000111100011000",
		b"11111110001010000111110110",
		b"11111110001011010111010010",
		b"11111110001100101010101001",
		b"11111110001110000001110111",
		b"11111110001111011100111001",
		b"11111110010000111011101010",
		b"11111110010010011110000111",
		b"11111110010100000100001011",
		b"11111110010101101101110010",
		b"11111110010111011010111000",
		b"11111110011001001011011000",
		b"11111110011010111111001101",
		b"11111110011100110110010011",
		b"11111110011110110000100101",
		b"11111110100000101101111111",
		b"11111110100010101110011010",
		b"11111110100100110001110010",
		b"11111110100110111000000010",
		b"11111110101001000001000100",
		b"11111110101011001100110011",
		b"11111110101101011011001010",
		b"11111110101111101100000011",
		b"11111110110001111111011000",
		b"11111110110100010101000100",
		b"11111110110110101101000001",
		b"11111110111001000111001010",
		b"11111110111011100011010111",
		b"11111110111110000001100100",
		b"11111111000000100001101011",
		b"11111111000011000011100100",
		b"11111111000101100111001100",
		b"11111111001000001100011010",
		b"11111111001010110011001001",
		b"11111111001101011011010011",
		b"11111111010000000100110010",
		b"11111111010010101111011111",
		b"11111111010101011011010100",
		b"11111111011000001000001010",
		b"11111111011010110101111100",
		b"11111111011101100100100011",
		b"11111111100000010011111001",
		b"11111111100011000011110111",
		b"11111111100101110100010111",
		b"11111111101000100101010011",
		b"11111111101011010110100100",
		b"11111111101110001000000100",
		b"11111111110000111001101100",
		b"11111111110011101011010110",
		b"11111111110110011100111101",
		b"11111111111001001110011001",
		b"11111111111011111111100100",
		b"11111111111110110000011000",
		b"00000000000001100000101111",
		b"00000000000100010000100011",
		b"00000000000110111111101101",
		b"00000000001001101110001000",
		b"00000000001100011011101101",
		b"00000000001111001000010110",
		b"00000000010001110011111110",
		b"00000000010100011110011110",
		b"00000000010111000111110001",
		b"00000000011001101111110000",
		b"00000000011100010110010111",
		b"00000000011110111011011111",
		b"00000000100001011111000011",
		b"00000000100100000000111101",
		b"00000000100110100001001000",
		b"00000000101000111111011110",
		b"00000000101011011011111011",
		b"00000000101101110110011001",
		b"00000000110000001110110010",
		b"00000000110010100101000011",
		b"00000000110100111001000101",
		b"00000000110111001010110100",
		b"00000000111001011010001100",
		b"00000000111011100111000111",
		b"00000000111101110001100001",
		b"00000000111111111001010110",
		b"00000001000001111110100001",
		b"00000001000100000000111110",
		b"00000001000110000000101001",
		b"00000001000111111101011101",
		b"00000001001001110111011000",
		b"00000001001011101110010101",
		b"00000001001101100010010000",
		b"00000001001111010011000110",
		b"00000001010001000000110100",
		b"00000001010010101011010101",
		b"00000001010100010010101000",
		b"00000001010101110110101000",
		b"00000001010111010111010011",
		b"00000001011000110100100111",
		b"00000001011010001110100000",
		b"00000001011011100100111011",
		b"00000001011100110111110111",
		b"00000001011110000111010001",
		b"00000001011111010011000111",
		b"00000001100000011011010111",
		b"00000001100001011111111110",
		b"00000001100010100000111100",
		b"00000001100011011110001111",
		b"00000001100100010111110100",
		b"00000001100101001101101011",
		b"00000001100101111111110011",
		b"00000001100110101110001010",
		b"00000001100111011000101111",
		b"00000001100111111111100010",
		b"00000001101000100010100010",
		b"00000001101001000001101110",
		b"00000001101001011101000110",
		b"00000001101001110100101010",
		b"00000001101010001000011001",
		b"00000001101010011000010100",
		b"00000001101010100100011010",
		b"00000001101010101100101101",
		b"00000001101010110001001011",
		b"00000001101010110001110111",
		b"00000001101010101110110000",
		b"00000001101010100111111000",
		b"00000001101010011101001110",
		b"00000001101010001110110110",
		b"00000001101001111100101110",
		b"00000001101001100110111010",
		b"00000001101001001101011010",
		b"00000001101000110000010000",
		b"00000001101000001111011101",
		b"00000001100111101011000100",
		b"00000001100111000011000111",
		b"00000001100110010111100111",
		b"00000001100101101000100110",
		b"00000001100100110110001000",
		b"00000001100100000000001110",
		b"00000001100011000110111011",
		b"00000001100010001010010001",
		b"00000001100001001010010100",
		b"00000001100000000111000111",
		b"00000001011111000000101011",
		b"00000001011101110111000101",
		b"00000001011100101010011000",
		b"00000001011011011010100110",
		b"00000001011010000111110011",
		b"00000001011000110010000011",
		b"00000001010111011001011010",
		b"00000001010101111101111010",
		b"00000001010100011111101001",
		b"00000001010010111110101001",
		b"00000001010001011010111110",
		b"00000001001111110100101101",
		b"00000001001110001011111010",
		b"00000001001100100000101000",
		b"00000001001010110010111101",
		b"00000001001001000010111100",
		b"00000001000111010000101010",
		b"00000001000101011100001011",
		b"00000001000011100101100101",
		b"00000001000001101100111010",
		b"00000000111111110010010001",
		b"00000000111101110101101110",
		b"00000000111011110111010101",
		b"00000000111001110111001100",
		b"00000000110111110101010111",
		b"00000000110101110001111011",
		b"00000000110011101100111110",
		b"00000000110001100110100100",
		b"00000000101111011110110001",
		b"00000000101101010101101101",
		b"00000000101011001011011010",
		b"00000000101000111111111111",
		b"00000000100110110011100001",
		b"00000000100100100110000100",
		b"00000000100010010111101111",
		b"00000000100000001000100110",
		b"00000000011101111000101110",
		b"00000000011011101000001101",
		b"00000000011001010111001000",
		b"00000000010111000101100100",
		b"00000000010100110011100110",
		b"00000000010010100001010100",
		b"00000000010000001110110100",
		b"00000000001101111100001001",
		b"00000000001011101001011010",
		b"00000000001001010110101011",
		b"00000000000111000100000010",
		b"00000000000100110001100100",
		b"00000000000010011111010110",
		b"00000000000000001101011110",
		b"11111111111101111100000000",
		b"11111111111011101011000001",
		b"11111111111001011010100111",
		b"11111111110111001010110111",
		b"11111111110100111011110101",
		b"11111111110010101101100110",
		b"11111111110000100000010000",
		b"11111111101110010011110111",
		b"11111111101100001000100000",
		b"11111111101001111110001111",
		b"11111111100111110101001010",
		b"11111111100101101101010110",
		b"11111111100011100110110101",
		b"11111111100001100001101110",
		b"11111111011111011110000101",
		b"11111111011101011011111101",
		b"11111111011011011011011100",
		b"11111111011001011100100110",
		b"11111111010111011111011110",
		b"11111111010101100100001001",
		b"11111111010011101010101011",
		b"11111111010001110011001000",
		b"11111111001111111101100100",
		b"11111111001110001010000010",
		b"11111111001100011000100111",
		b"11111111001010101001010101",
		b"11111111001000111100010001",
		b"11111111000111010001011110",
		b"11111111000101101000111111",
		b"11111111000100000010110111",
		b"11111111000010011111001011",
		b"11111111000000111101111100",
		b"11111110111111011111001101",
		b"11111110111110000011000011",
		b"11111110111100101001011111",
		b"11111110111011010010100100",
		b"11111110111001111110010100",
		b"11111110111000101100110011",
		b"11111110110111011110000011",
		b"11111110110110010010000101",
		b"11111110110101001000111100",
		b"11111110110100000010101011",
		b"11111110110010111111010010",
		b"11111110110001111110110101",
		b"11111110110001000001010100",
		b"11111110110000000110110001",
		b"11111110101111001111001110",
		b"11111110101110011010101100",
		b"11111110101101101001001100",
		b"11111110101100111010110001",
		b"11111110101100001111011010",
		b"11111110101011100111001000",
		b"11111110101011000001111101",
		b"11111110101010011111111010",
		b"11111110101010000000111110",
		b"11111110101001100101001011",
		b"11111110101001001100100001",
		b"11111110101000110110111111",
		b"11111110101000100100100111",
		b"11111110101000010101011000",
		b"11111110101000001001010011",
		b"11111110101000000000010110",
		b"11111110100111111010100011",
		b"11111110100111110111110111",
		b"11111110100111111000010100",
		b"11111110100111111011111000",
		b"11111110101000000010100011",
		b"11111110101000001100010100",
		b"11111110101000011001001001",
		b"11111110101000101001000011",
		b"11111110101000111011111111",
		b"11111110101001010001111101",
		b"11111110101001101010111010",
		b"11111110101010000110110111",
		b"11111110101010100101110000",
		b"11111110101011000111100110",
		b"11111110101011101100010100",
		b"11111110101100010011111011",
		b"11111110101100111110011000",
		b"11111110101101101011101001",
		b"11111110101110011011101011",
		b"11111110101111001110011101",
		b"11111110110000000011111101",
		b"11111110110000111100000111",
		b"11111110110001110110111001",
		b"11111110110010110100010010",
		b"11111110110011110100001101",
		b"11111110110100110110101001",
		b"11111110110101111011100011",
		b"11111110110111000010110111",
		b"11111110111000001100100010",
		b"11111110111001011000100011",
		b"11111110111010100110110101",
		b"11111110111011110111010101",
		b"11111110111101001010000000",
		b"11111110111110011110110011",
		b"11111110111111110101101011",
		b"11111111000001001110100011",
		b"11111111000010101001011000",
		b"11111111000100000110001000",
		b"11111111000101100100101101",
		b"11111111000111000101000101",
		b"11111111001000100111001011",
		b"11111111001010001010111100",
		b"11111111001011110000010101",
		b"11111111001101010111010000",
		b"11111111001110111111101011",
		b"11111111010000101001100000",
		b"11111111010010010100101101",
		b"11111111010100000001001110",
		b"11111111010101101110111101",
		b"11111111010111011101110111",
		b"11111111011001001101111000",
		b"11111111011010111110111100",
		b"11111111011100110000111110",
		b"11111111011110100011111010",
		b"11111111100000010111101100",
		b"11111111100010001100010000",
		b"11111111100100000001100010",
		b"11111111100101110111011101",
		b"11111111100111101101111100",
		b"11111111101001100100111101",
		b"11111111101011011100011001",
		b"11111111101101010100001110",
		b"11111111101111001100010110",
		b"11111111110001000100101101",
		b"11111111110010111101010000",
		b"11111111110100110101111001",
		b"11111111110110101110100101",
		b"11111111111000100111001111",
		b"11111111111010011111110011",
		b"11111111111100011000001101",
		b"11111111111110010000011000",
		b"00000000000000001000010001",
		b"00000000000001111111110010",
		b"00000000000011110110111001",
		b"00000000000101101101100000",
		b"00000000000111100011100100",
		b"00000000001001011001000001",
		b"00000000001011001101110010",
		b"00000000001101000001110100",
		b"00000000001110110101000011",
		b"00000000010000100111011010",
		b"00000000010010011000110110",
		b"00000000010100001001010011",
		b"00000000010101111000101110",
		b"00000000010111100111000010",
		b"00000000011001010100001011",
		b"00000000011011000000000111",
		b"00000000011100101010110010",
		b"00000000011110010100000111",
		b"00000000011111111100000100",
		b"00000000100001100010100110",
		b"00000000100011000111101000",
		b"00000000100100101011000111",
		b"00000000100110001101000001",
		b"00000000100111101101010010",
		b"00000000101001001011111000",
		b"00000000101010101000101110",
		b"00000000101100000011110010",
		b"00000000101101011101000010",
		b"00000000101110110100011010",
		b"00000000110000001001111000",
		b"00000000110001011101011000",
		b"00000000110010101110111010",
		b"00000000110011111110011001",
		b"00000000110101001011110100",
		b"00000000110110010111000111",
		b"00000000110111100000010010",
		b"00000000111000100111010010",
		b"00000000111001101100000100",
		b"00000000111010101110100111",
		b"00000000111011101110111001",
		b"00000000111100101100111000",
		b"00000000111101101000100010",
		b"00000000111110100001110101",
		b"00000000111111011000110000",
		b"00000001000000001101010010",
		b"00000001000000111111011001",
		b"00000001000001101111000011",
		b"00000001000010011100010001",
		b"00000001000011000110111111",
		b"00000001000011101111001110",
		b"00000001000100010100111100",
		b"00000001000100111000001001",
		b"00000001000101011000110100",
		b"00000001000101110110111100",
		b"00000001000110010010100000",
		b"00000001000110101011100001",
		b"00000001000111000001111101",
		b"00000001000111010101110101",
		b"00000001000111100111001000",
		b"00000001000111110101110110",
		b"00000001001000000001111111",
		b"00000001001000001011100011",
		b"00000001001000010010100011",
		b"00000001001000010110111110",
		b"00000001001000011000110100",
		b"00000001001000011000001000",
		b"00000001001000010100111000",
		b"00000001001000001111000101",
		b"00000001001000000110110001",
		b"00000001000111111011111011",
		b"00000001000111101110100110",
		b"00000001000111011110110001",
		b"00000001000111001100011101",
		b"00000001000110110111101101",
		b"00000001000110100000100001",
		b"00000001000110000110111010",
		b"00000001000101101010111010",
		b"00000001000101001100100010",
		b"00000001000100101011110011",
		b"00000001000100001000110001",
		b"00000001000011100011011011",
		b"00000001000010111011110100",
		b"00000001000010010001111101",
		b"00000001000001100101111001",
		b"00000001000000110111101010",
		b"00000001000000000111010001",
		b"00000000111111010100110001",
		b"00000000111110100000001100",
		b"00000000111101101001100100",
		b"00000000111100110000111011",
		b"00000000111011110110010100",
		b"00000000111010111001110010",
		b"00000000111001111011010110",
		b"00000000111000111011000100",
		b"00000000110111111000111101",
		b"00000000110110110101000110",
		b"00000000110101101111100000",
		b"00000000110100101000001110",
		b"00000000110011011111010011",
		b"00000000110010010100110010",
		b"00000000110001001000101101",
		b"00000000101111111011001001",
		b"00000000101110101100001000",
		b"00000000101101011011101100",
		b"00000000101100001001111010",
		b"00000000101010110110110100",
		b"00000000101001100010011101",
		b"00000000101000001100111001",
		b"00000000100110110110001011",
		b"00000000100101011110010110",
		b"00000000100100000101011101",
		b"00000000100010101011100101",
		b"00000000100001010000101111",
		b"00000000011111110101000000",
		b"00000000011110011000011011",
		b"00000000011100111011000011",
		b"00000000011011011100111101",
		b"00000000011001111110001010",
		b"00000000011000011110101111",
		b"00000000010110111110110000",
		b"00000000010101011110001111",
		b"00000000010011111101010001",
		b"00000000010010011011111000",
		b"00000000010000111010001001",
		b"00000000001111011000000110",
		b"00000000001101110101110100",
		b"00000000001100010011010110",
		b"00000000001010110000101111",
		b"00000000001001001110000011",
		b"00000000000111101011010101",
		b"00000000000110001000101001",
		b"00000000000100100110000010",
		b"00000000000011000011100100",
		b"00000000000001100001010010",
		b"11111111111111111111010000",
		b"11111111111110011101100001",
		b"11111111111100111100001000",
		b"11111111111011011011001001",
		b"11111111111001111010100111",
		b"11111111111000011010100110",
		b"11111111110110111011001000",
		b"11111111110101011100010010",
		b"11111111110011111110000101",
		b"11111111110010100000100110",
		b"11111111110001000011110111",
		b"11111111101111100111111100",
		b"11111111101110001100111000",
		b"11111111101100110010101110",
		b"11111111101011011001100000",
		b"11111111101010000001010010",
		b"11111111101000101010000111",
		b"11111111100111010100000001",
		b"11111111100101111111000100",
		b"11111111100100101011010001",
		b"11111111100011011000101101",
		b"11111111100010000111011001",
		b"11111111100000110111011000",
		b"11111111011111101000101101",
		b"11111111011110011011011010",
		b"11111111011101001111100001",
		b"11111111011100000101000110",
		b"11111111011010111100001010",
		b"11111111011001110100110000",
		b"11111111011000101110111001",
		b"11111111010111101010101000",
		b"11111111010110101000000000",
		b"11111111010101100111000010",
		b"11111111010100100111101111",
		b"11111111010011101010001011",
		b"11111111010010101110010111",
		b"11111111010001110100010100",
		b"11111111010000111100000100",
		b"11111111010000000101101001",
		b"11111111001111010001000101",
		b"11111111001110011110011001",
		b"11111111001101101101100110",
		b"11111111001100111110101101",
		b"11111111001100010001110001",
		b"11111111001011100110110010",
		b"11111111001010111101110001",
		b"11111111001010010110101111",
		b"11111111001001110001101110",
		b"11111111001001001110101110",
		b"11111111001000101101110000",
		b"11111111001000001110110101",
		b"11111111000111110001111101",
		b"11111111000111010111001001",
		b"11111111000110111110011011",
		b"11111111000110100111110001",
		b"11111111000110010011001100",
		b"11111111000110000000101110",
		b"11111111000101110000010101",
		b"11111111000101100010000011",
		b"11111111000101010101110111",
		b"11111111000101001011110010",
		b"11111111000101000011110010",
		b"11111111000100111101111001",
		b"11111111000100111010000101",
		b"11111111000100111000011000",
		b"11111111000100111000101111",
		b"11111111000100111011001011",
		b"11111111000100111111101100",
		b"11111111000101000110010000",
		b"11111111000101001110111000",
		b"11111111000101011001100010",
		b"11111111000101100110001101",
		b"11111111000101110100111010",
		b"11111111000110000101100110",
		b"11111111000110011000010001",
		b"11111111000110101100111010",
		b"11111111000111000011100000",
		b"11111111000111011100000001",
		b"11111111000111110110011101",
		b"11111111001000010010110001",
		b"11111111001000110000111101",
		b"11111111001001010001000000",
		b"11111111001001110010110111",
		b"11111111001010010110100001",
		b"11111111001010111011111101",
		b"11111111001011100011001000",
		b"11111111001100001100000010",
		b"11111111001100110110101000",
		b"11111111001101100010111000",
		b"11111111001110010000110001",
		b"11111111001111000000010001",
		b"11111111001111110001010101",
		b"11111111010000100011111100",
		b"11111111010001011000000100",
		b"11111111010010001101101010",
		b"11111111010011000100101100",
		b"11111111010011111101001001",
		b"11111111010100110110111101",
		b"11111111010101110010000111",
		b"11111111010110101110100011",
		b"11111111010111101100010001",
		b"11111111011000101011001100",
		b"11111111011001101011010100",
		b"11111111011010101100100101",
		b"11111111011011101110111101",
		b"11111111011100110010011001",
		b"11111111011101110110110110",
		b"11111111011110111100010011",
		b"11111111100000000010101100",
		b"11111111100001001001111111",
		b"11111111100010010010001001",
		b"11111111100011011011001000",
		b"11111111100100100100111000",
		b"11111111100101101111010111",
		b"11111111100110111010100010",
		b"11111111101000000110010111",
		b"11111111101001010010110010",
		b"11111111101010011111110001",
		b"11111111101011101101010001",
		b"11111111101100111011001111",
		b"11111111101110001001101000",
		b"11111111101111011000011010",
		b"11111111110000100111100010",
		b"11111111110001110110111100",
		b"11111111110011000110100110",
		b"11111111110100010110011101",
		b"11111111110101100110011110",
		b"11111111110110110110100111",
		b"11111111111000000110110100",
		b"11111111111001010111000011",
		b"11111111111010100111010001",
		b"11111111111011110111011011",
		b"11111111111101000111011110",
		b"11111111111110010111011000",
		b"11111111111111100111000110",
		b"00000000000000110110100100",
		b"00000000000010000101110001",
		b"00000000000011010100101001",
		b"00000000000100100011001001",
		b"00000000000101110001010000",
		b"00000000000110111110111011",
		b"00000000001000001100000110",
		b"00000000001001011000101111",
		b"00000000001010100100110100",
		b"00000000001011110000010010",
		b"00000000001100111011000111",
		b"00000000001110000101001111",
		b"00000000001111001110101001",
		b"00000000010000010111010010",
		b"00000000010001011111001000",
		b"00000000010010100110001001",
		b"00000000010011101100010001",
		b"00000000010100110001011111",
		b"00000000010101110101110001",
		b"00000000010110111001000100",
		b"00000000010111111011010110",
		b"00000000011000111100100110",
		b"00000000011001111100110000",
		b"00000000011010111011110011",
		b"00000000011011111001101101",
		b"00000000011100110110011100",
		b"00000000011101110001111110",
		b"00000000011110101100010010",
		b"00000000011111100101010101",
		b"00000000100000011101000101",
		b"00000000100001010011100010",
		b"00000000100010001000101001",
		b"00000000100010111100011001",
		b"00000000100011101110110000",
		b"00000000100100011111101101",
		b"00000000100101001111001110",
		b"00000000100101111101010010",
		b"00000000100110101001111000",
		b"00000000100111010100111110",
		b"00000000100111111110100100",
		b"00000000101000100110100111",
		b"00000000101001001101001000",
		b"00000000101001110010000100",
		b"00000000101010010101011011",
		b"00000000101010110111001101",
		b"00000000101011010111010111",
		b"00000000101011110101111010",
		b"00000000101100010010110100",
		b"00000000101100101110000101",
		b"00000000101101000111101101",
		b"00000000101101011111101010",
		b"00000000101101110101111101",
		b"00000000101110001010100100",
		b"00000000101110011101100000",
		b"00000000101110101110110000",
		b"00000000101110111110010100",
		b"00000000101111001100001011",
		b"00000000101111011000010110",
		b"00000000101111100010110100",
		b"00000000101111101011100110",
		b"00000000101111110010101011",
		b"00000000101111111000000100",
		b"00000000101111111011110001",
		b"00000000101111111101110001",
		b"00000000101111111110000110",
		b"00000000101111111100101111",
		b"00000000101111111001101101",
		b"00000000101111110101000000",
		b"00000000101111101110101001",
		b"00000000101111100110101001",
		b"00000000101111011101000000",
		b"00000000101111010001101110",
		b"00000000101111000100110101",
		b"00000000101110110110010110",
		b"00000000101110100110010000",
		b"00000000101110010100100101",
		b"00000000101110000001010110",
		b"00000000101101101100100101",
		b"00000000101101010110010001",
		b"00000000101100111110011100",
		b"00000000101100100101000111",
		b"00000000101100001010010100",
		b"00000000101011101110000011",
		b"00000000101011010000010111",
		b"00000000101010110001001111",
		b"00000000101010010000101111",
		b"00000000101001101110110110",
		b"00000000101001001011100111",
		b"00000000101000100111000011",
		b"00000000101000000001001100",
		b"00000000100111011010000010",
		b"00000000100110110001101001",
		b"00000000100110001000000001",
		b"00000000100101011101001100",
		b"00000000100100110001001101",
		b"00000000100100000100000100",
		b"00000000100011010101110100",
		b"00000000100010100110011110",
		b"00000000100001110110000100",
		b"00000000100001000100101001",
		b"00000000100000010010001101",
		b"00000000011111011110110100",
		b"00000000011110101010011111",
		b"00000000011101110101010001",
		b"00000000011100111111001010",
		b"00000000011100001000001110",
		b"00000000011011010000011110",
		b"00000000011010010111111100",
		b"00000000011001011110101011",
		b"00000000011000100100101101",
		b"00000000010111101010000100",
		b"00000000010110101110110010",
		b"00000000010101110010111010",
		b"00000000010100110110011101",
		b"00000000010011111001011110",
		b"00000000010010111011111111",
		b"00000000010001111110000010",
		b"00000000010000111111101001",
		b"00000000010000000000111000",
		b"00000000001111000001110000",
		b"00000000001110000010010011",
		b"00000000001101000010100100",
		b"00000000001100000010100101",
		b"00000000001011000010011000",
		b"00000000001010000001111111",
		b"00000000001001000001011110",
		b"00000000001000000000110101",
		b"00000000000111000000001000",
		b"00000000000101111111011001",
		b"00000000000100111110101010",
		b"00000000000011111101111101",
		b"00000000000010111101010100",
		b"00000000000001111100110010",
		b"00000000000000111100011001",
		b"11111111111111111100001100",
		b"11111111111110111100001011",
		b"11111111111101111100011011",
		b"11111111111100111100111100",
		b"11111111111011111101110001",
		b"11111111111010111110111100",
		b"11111111111010000000011111",
		b"11111111111001000010011100",
		b"11111111111000000100110110",
		b"11111111110111000111101110",
		b"11111111110110001011000111",
		b"11111111110101001111000011",
		b"11111111110100010011100010",
		b"11111111110011011000101000",
		b"11111111110010011110010111",
		b"11111111110001100100110000",
		b"11111111110000101011110101",
		b"11111111101111110011101000",
		b"11111111101110111100001010",
		b"11111111101110000101011111",
		b"11111111101101001111100110",
		b"11111111101100011010100011",
		b"11111111101011100110010110",
		b"11111111101010110011000010",
		b"11111111101010000000101000",
		b"11111111101001001111001001",
		b"11111111101000011110100111",
		b"11111111100111101111000100",
		b"11111111100111000000100001",
		b"11111111100110010011000000",
		b"11111111100101100110100001",
		b"11111111100100111011000110",
		b"11111111100100010000110001",
		b"11111111100011100111100010",
		b"11111111100010111111011100",
		b"11111111100010011000011110",
		b"11111111100001110010101011",
		b"11111111100001001110000011",
		b"11111111100000101010100111",
		b"11111111100000001000011000",
		b"11111111011111100111011000",
		b"11111111011111000111100110",
		b"11111111011110101001000101",
		b"11111111011110001011110101",
		b"11111111011101101111110110",
		b"11111111011101010101001001",
		b"11111111011100111011101111",
		b"11111111011100100011101000",
		b"11111111011100001100110110",
		b"11111111011011110111011000",
		b"11111111011011100011001111",
		b"11111111011011010000011100",
		b"11111111011010111110111110",
		b"11111111011010101110110111",
		b"11111111011010100000000110",
		b"11111111011010010010101100",
		b"11111111011010000110101001",
		b"11111111011001111011111100",
		b"11111111011001110010100111",
		b"11111111011001101010101001",
		b"11111111011001100100000010",
		b"11111111011001011110110010",
		b"11111111011001011010111000",
		b"11111111011001011000010110",
		b"11111111011001010111001010",
		b"11111111011001010111010101",
		b"11111111011001011000110110",
		b"11111111011001011011101100",
		b"11111111011001011111111000",
		b"11111111011001100101011000",
		b"11111111011001101100001101",
		b"11111111011001110100010110",
		b"11111111011001111101110010",
		b"11111111011010001000100001",
		b"11111111011010010100100010",
		b"11111111011010100001110100",
		b"11111111011010110000011000",
		b"11111111011011000000001010",
		b"11111111011011010001001100",
		b"11111111011011100011011101",
		b"11111111011011110110111010",
		b"11111111011100001011100100",
		b"11111111011100100001011001",
		b"11111111011100111000011001",
		b"11111111011101010000100010",
		b"11111111011101101001110011",
		b"11111111011110000100001100",
		b"11111111011110011111101010",
		b"11111111011110111100001101",
		b"11111111011111011001110100",
		b"11111111011111111000011101",
		b"11111111100000011000000111",
		b"11111111100000111000110001",
		b"11111111100001011010011001",
		b"11111111100001111100111110",
		b"11111111100010100000011111",
		b"11111111100011000100111010",
		b"11111111100011101010001101",
		b"11111111100100010000011000",
		b"11111111100100110111011000",
		b"11111111100101011111001100",
		b"11111111100110000111110011",
		b"11111111100110110001001011",
		b"11111111100111011011010010",
		b"11111111101000000110000111",
		b"11111111101000110001101000",
		b"11111111101001011101110100",
		b"11111111101010001010101000",
		b"11111111101010111000000100",
		b"11111111101011100110000100",
		b"11111111101100010100101001",
		b"11111111101101000011101111",
		b"11111111101101110011010101",
		b"11111111101110100011011010",
		b"11111111101111010011111011",
		b"11111111110000000100110111",
		b"11111111110000110110001100",
		b"11111111110001100111111000",
		b"11111111110010011001111010",
		b"11111111110011001100001111",
		b"11111111110011111110110110",
		b"11111111110100110001101101",
		b"11111111110101100100110010",
		b"11111111110110011000000100",
		b"11111111110111001011100000",
		b"11111111110111111111000100",
		b"11111111111000110010110000",
		b"11111111111001100110100000",
		b"11111111111010011010010011",
		b"11111111111011001110001000",
		b"11111111111100000001111101",
		b"11111111111100110101101111",
		b"11111111111101101001011101",
		b"11111111111110011101000110",
		b"11111111111111010000100110",
		b"00000000000000000011111110",
		b"00000000000000110111001010",
		b"00000000000001101010001010",
		b"00000000000010011100111011",
		b"00000000000011001111011011",
		b"00000000000100000001101010",
		b"00000000000100110011100101",
		b"00000000000101100101001011",
		b"00000000000110010110011001",
		b"00000000000111000111001111",
		b"00000000000111110111101011",
		b"00000000001000100111101011",
		b"00000000001001010111001101",
		b"00000000001010000110010000",
		b"00000000001010110100110011",
		b"00000000001011100010110100",
		b"00000000001100010000010010",
		b"00000000001100111101001010",
		b"00000000001101101001011100",
		b"00000000001110010101000111",
		b"00000000001111000000001000",
		b"00000000001111101010011110",
		b"00000000010000010100001001",
		b"00000000010000111101000111",
		b"00000000010001100101010110",
		b"00000000010010001100110101",
		b"00000000010010110011100100",
		b"00000000010011011001100000",
		b"00000000010011111110101010",
		b"00000000010100100010111111",
		b"00000000010101000110011110",
		b"00000000010101101001001000",
		b"00000000010110001010111001",
		b"00000000010110101011110010",
		b"00000000010111001011110010",
		b"00000000010111101010111000",
		b"00000000011000001001000010",
		b"00000000011000100110010000",
		b"00000000011001000010100010",
		b"00000000011001011101110101",
		b"00000000011001111000001011",
		b"00000000011010010001100001",
		b"00000000011010101001110111",
		b"00000000011011000001001110",
		b"00000000011011010111100011",
		b"00000000011011101100110111",
		b"00000000011100000001001000",
		b"00000000011100010100011000",
		b"00000000011100100110100100",
		b"00000000011100110111101101",
		b"00000000011101000111110010",
		b"00000000011101010110110011",
		b"00000000011101100100110000",
		b"00000000011101110001101000",
		b"00000000011101111101011100",
		b"00000000011110001000001010",
		b"00000000011110010001110100",
		b"00000000011110011010011000",
		b"00000000011110100001110111",
		b"00000000011110101000010001",
		b"00000000011110101101100101",
		b"00000000011110110001110100",
		b"00000000011110110100111111",
		b"00000000011110110111000100",
		b"00000000011110111000000100",
		b"00000000011110111000000000",
		b"00000000011110110110110111",
		b"00000000011110110100101010",
		b"00000000011110110001011010",
		b"00000000011110101101000110",
		b"00000000011110100111101111",
		b"00000000011110100001010101",
		b"00000000011110011001111001",
		b"00000000011110010001011011",
		b"00000000011110000111111100",
		b"00000000011101111101011101",
		b"00000000011101110001111101",
		b"00000000011101100101011110",
		b"00000000011101011000000000",
		b"00000000011101001001100100",
		b"00000000011100111010001011",
		b"00000000011100101001110101",
		b"00000000011100011000100011",
		b"00000000011100000110010111",
		b"00000000011011110011001111",
		b"00000000011011011111001111",
		b"00000000011011001010010110",
		b"00000000011010110100100110",
		b"00000000011010011101111110",
		b"00000000011010000110100010",
		b"00000000011001101110010000",
		b"00000000011001010101001011",
		b"00000000011000111011010100",
		b"00000000011000100000101011",
		b"00000000011000000101010001",
		b"00000000010111101001001000",
		b"00000000010111001100010010",
		b"00000000010110101110101110",
		b"00000000010110010000011110",
		b"00000000010101110001100100",
		b"00000000010101010010000000",
		b"00000000010100110001110100",
		b"00000000010100010001000001",
		b"00000000010011101111101001",
		b"00000000010011001101101100",
		b"00000000010010101011001100",
		b"00000000010010001000001011",
		b"00000000010001100100101001",
		b"00000000010001000000101000",
		b"00000000010000011100001001",
		b"00000000001111110111001110",
		b"00000000001111010001111000",
		b"00000000001110101100001000",
		b"00000000001110000110000000",
		b"00000000001101011111100010",
		b"00000000001100111000101110",
		b"00000000001100010001100110",
		b"00000000001011101010001011",
		b"00000000001011000010100000",
		b"00000000001010011010100101",
		b"00000000001001110010011011",
		b"00000000001001001010000101",
		b"00000000001000100001100011",
		b"00000000000111111000111000",
		b"00000000000111010000000100",
		b"00000000000110100111001001",
		b"00000000000101111110001000",
		b"00000000000101010101000100",
		b"00000000000100101011111100",
		b"00000000000100000010110011",
		b"00000000000011011001101011",
		b"00000000000010110000100100",
		b"00000000000010000111011111",
		b"00000000000001011110100000",
		b"00000000000000110101100110",
		b"00000000000000001100110011",
		b"11111111111111100100001001",
		b"11111111111110111011101001",
		b"11111111111110010011010100",
		b"11111111111101101011001011",
		b"11111111111101000011010001",
		b"11111111111100011011100110",
		b"11111111111011110100001100",
		b"11111111111011001101000011",
		b"11111111111010100110001110",
		b"11111111111001111111101110",
		b"11111111111001011001100011",
		b"11111111111000110011101111",
		b"11111111111000001110010011",
		b"11111111110111101001010001",
		b"11111111110111000100101010",
		b"11111111110110100000011110",
		b"11111111110101111100101111",
		b"11111111110101011001011111",
		b"11111111110100110110101101",
		b"11111111110100010100011100",
		b"11111111110011110010101100",
		b"11111111110011010001011111",
		b"11111111110010110000110101",
		b"11111111110010010000110000",
		b"11111111110001110001010000",
		b"11111111110001010010010110",
		b"11111111110000110100000100",
		b"11111111110000010110011001",
		b"11111111101111111001011000",
		b"11111111101111011101000001",
		b"11111111101111000001010101",
		b"11111111101110100110010100",
		b"11111111101110001100000000",
		b"11111111101101110010011001",
		b"11111111101101011001011111",
		b"11111111101101000001010100",
		b"11111111101100101001111001",
		b"11111111101100010011001101",
		b"11111111101011111101010010",
		b"11111111101011101000000111",
		b"11111111101011010011101111",
		b"11111111101011000000001000",
		b"11111111101010101101010100",
		b"11111111101010011011010011",
		b"11111111101010001010000110",
		b"11111111101001111001101101",
		b"11111111101001101010001000",
		b"11111111101001011011011000",
		b"11111111101001001101011100",
		b"11111111101001000000010111",
		b"11111111101000110100000110",
		b"11111111101000101000101100",
		b"11111111101000011110000111",
		b"11111111101000010100011001",
		b"11111111101000001011100001",
		b"11111111101000000011011111",
		b"11111111100111111100010100",
		b"11111111100111110101111111",
		b"11111111100111110000100001",
		b"11111111100111101011111010",
		b"11111111100111101000001001",
		b"11111111100111100101001111",
		b"11111111100111100011001011",
		b"11111111100111100001111110",
		b"11111111100111100001100110",
		b"11111111100111100010000100",
		b"11111111100111100011011001",
		b"11111111100111100101100010",
		b"11111111100111101000100001",
		b"11111111100111101100010101",
		b"11111111100111110000111110",
		b"11111111100111110110011010",
		b"11111111100111111100101011",
		b"11111111101000000011101111",
		b"11111111101000001011100111",
		b"11111111101000010100010001",
		b"11111111101000011101101101",
		b"11111111101000100111111010",
		b"11111111101000110010111001",
		b"11111111101000111110101001",
		b"11111111101001001011001000",
		b"11111111101001011000010111",
		b"11111111101001100110010100",
		b"11111111101001110101000000",
		b"11111111101010000100011001",
		b"11111111101010010100011111",
		b"11111111101010100101010001",
		b"11111111101010110110101110",
		b"11111111101011001000110110",
		b"11111111101011011011100111",
		b"11111111101011101111000010",
		b"11111111101100000011000100",
		b"11111111101100010111101110",
		b"11111111101100101100111111",
		b"11111111101101000010110101",
		b"11111111101101011001010000",
		b"11111111101101110000001110",
		b"11111111101110000111110000",
		b"11111111101110011111110011",
		b"11111111101110111000011000",
		b"11111111101111010001011100",
		b"11111111101111101011000000",
		b"11111111110000000101000010",
		b"11111111110000011111100001",
		b"11111111110000111010011100",
		b"11111111110001010101110010",
		b"11111111110001110001100010",
		b"11111111110010001101101011",
		b"11111111110010101010001100",
		b"11111111110011000111000011",
		b"11111111110011100100010001",
		b"11111111110100000001110011",
		b"11111111110100011111101001",
		b"11111111110100111101110001",
		b"11111111110101011100001011",
		b"11111111110101111010110101",
		b"11111111110110011001101110",
		b"11111111110110111000110110",
		b"11111111110111011000001010",
		b"11111111110111110111101010",
		b"11111111111000010111010101",
		b"11111111111000110111001001",
		b"11111111111001010111000110",
		b"11111111111001110111001010",
		b"11111111111010010111010100",
		b"11111111111010110111100100",
		b"11111111111011010111110111",
		b"11111111111011111000001101",
		b"11111111111100011000100101",
		b"11111111111100111000111110",
		b"11111111111101011001010110",
		b"11111111111101111001101100",
		b"11111111111110011010000000",
		b"11111111111110111010001111",
		b"11111111111111011010011010",
		b"11111111111111111010011111",
		b"00000000000000011010011101",
		b"00000000000000111010010010",
		b"00000000000001011001111110",
		b"00000000000001111001100000",
		b"00000000000010011000110111",
		b"00000000000010111000000001",
		b"00000000000011010110111110",
		b"00000000000011110101101101",
		b"00000000000100010100001100",
		b"00000000000100110010011011",
		b"00000000000101010000011000",
		b"00000000000101101110000011",
		b"00000000000110001011011011",
		b"00000000000110101000011111",
		b"00000000000111000101001101",
		b"00000000000111100001100101",
		b"00000000000111111101100111",
		b"00000000001000011001010000",
		b"00000000001000110100100001",
		b"00000000001001001111011001",
		b"00000000001001101001110110",
		b"00000000001010000011110111",
		b"00000000001010011101011101",
		b"00000000001010110110100110",
		b"00000000001011001111010010",
		b"00000000001011100111100000",
		b"00000000001011111111001110",
		b"00000000001100010110011101",
		b"00000000001100101101001011",
		b"00000000001101000011011001",
		b"00000000001101011001000101",
		b"00000000001101101110001110",
		b"00000000001110000010110101",
		b"00000000001110010110111000",
		b"00000000001110101010011000",
		b"00000000001110111101010010",
		b"00000000001111001111101000",
		b"00000000001111100001011000",
		b"00000000001111110010100010",
		b"00000000010000000011000110",
		b"00000000010000010011000011",
		b"00000000010000100010011001",
		b"00000000010000110001000110",
		b"00000000010000111111001100",
		b"00000000010001001100101010",
		b"00000000010001011001011111",
		b"00000000010001100101101010",
		b"00000000010001110001001101",
		b"00000000010001111100000110",
		b"00000000010010000110010101",
		b"00000000010010001111111011",
		b"00000000010010011000110110",
		b"00000000010010100001001000",
		b"00000000010010101000101110",
		b"00000000010010101111101011",
		b"00000000010010110101111100",
		b"00000000010010111011100100",
		b"00000000010011000000100000",
		b"00000000010011000100110010",
		b"00000000010011001000011001",
		b"00000000010011001011010110",
		b"00000000010011001101101000",
		b"00000000010011001111001111",
		b"00000000010011010000001100",
		b"00000000010011010000011111",
		b"00000000010011010000001000",
		b"00000000010011001111000111",
		b"00000000010011001101011100",
		b"00000000010011001011000111",
		b"00000000010011001000001010",
		b"00000000010011000100100011",
		b"00000000010011000000010011",
		b"00000000010010111011011011",
		b"00000000010010110101111010",
		b"00000000010010101111110010",
		b"00000000010010101001000010",
		b"00000000010010100001101011",
		b"00000000010010011001101101",
		b"00000000010010010001001001",
		b"00000000010010001000000000",
		b"00000000010001111110010000",
		b"00000000010001110011111100",
		b"00000000010001101001000011",
		b"00000000010001011101100110",
		b"00000000010001010001100110",
		b"00000000010001000101000011",
		b"00000000010000110111111101",
		b"00000000010000101010010110",
		b"00000000010000011100001110",
		b"00000000010000001101100100",
		b"00000000001111111110011011",
		b"00000000001111101110110011",
		b"00000000001111011110101100",
		b"00000000001111001110000111",
		b"00000000001110111101000100",
		b"00000000001110101011100101",
		b"00000000001110011001101010",
		b"00000000001110000111010011",
		b"00000000001101110100100010",
		b"00000000001101100001011000",
		b"00000000001101001101110100",
		b"00000000001100111001111000",
		b"00000000001100100101100100",
		b"00000000001100010000111010",
		b"00000000001011111011111001",
		b"00000000001011100110100100",
		b"00000000001011010000111010",
		b"00000000001010111010111101",
		b"00000000001010100100101100",
		b"00000000001010001110001010",
		b"00000000001001110111010111",
		b"00000000001001100000010100",
		b"00000000001001001001000001",
		b"00000000001000110001100000",
		b"00000000001000011001110001",
		b"00000000001000000001110101",
		b"00000000000111101001101110",
		b"00000000000111010001011011",
		b"00000000000110111000111110",
		b"00000000000110100000011000",
		b"00000000000110000111101001",
		b"00000000000101101110110010",
		b"00000000000101010101110101",
		b"00000000000100111100110010",
		b"00000000000100100011101010",
		b"00000000000100001010011110",
		b"00000000000011110001001111",
		b"00000000000011010111111101",
		b"00000000000010111110101010",
		b"00000000000010100101010110",
		b"00000000000010001100000010",
		b"00000000000001110010101111",
		b"00000000000001011001011111",
		b"00000000000001000000010001",
		b"00000000000000100111000111",
		b"00000000000000001110000001",
		b"11111111111111110101000000",
		b"11111111111111011100000110",
		b"11111111111111000011010011",
		b"11111111111110101010100111",
		b"11111111111110010010000100",
		b"11111111111101111001101011",
		b"11111111111101100001011011",
		b"11111111111101001001010111",
		b"11111111111100110001011111",
		b"11111111111100011001110010",
		b"11111111111100000010010100",
		b"11111111111011101011000011",
		b"11111111111011010100000001",
		b"11111111111010111101001110",
		b"11111111111010100110101100",
		b"11111111111010010000011011",
		b"11111111111001111010011011",
		b"11111111111001100100101110",
		b"11111111111001001111010011",
		b"11111111111000111010001100",
		b"11111111111000100101011010",
		b"11111111111000010000111100",
		b"11111111110111111100110100",
		b"11111111110111101001000010",
		b"11111111110111010101100110",
		b"11111111110111000010100010",
		b"11111111110110101111110110",
		b"11111111110110011101100010",
		b"11111111110110001011100111",
		b"11111111110101111010000110",
		b"11111111110101101000111111",
		b"11111111110101011000010001",
		b"11111111110101000111111111",
		b"11111111110100111000001000",
		b"11111111110100101000101101",
		b"11111111110100011001101111",
		b"11111111110100001011001100",
		b"11111111110011111101000111",
		b"11111111110011101111011111",
		b"11111111110011100010010101",
		b"11111111110011010101101001",
		b"11111111110011001001011011",
		b"11111111110010111101101100",
		b"11111111110010110010011100",
		b"11111111110010100111101011",
		b"11111111110010011101011010",
		b"11111111110010010011101000",
		b"11111111110010001010010110",
		b"11111111110010000001100101",
		b"11111111110001111001010011",
		b"11111111110001110001100010",
		b"11111111110001101010010010",
		b"11111111110001100011100011",
		b"11111111110001011101010100",
		b"11111111110001010111100110",
		b"11111111110001010010011001",
		b"11111111110001001101101110",
		b"11111111110001001001100011",
		b"11111111110001000101111010",
		b"11111111110001000010110001",
		b"11111111110001000000001010",
		b"11111111110000111110000100",
		b"11111111110000111100011110",
		b"11111111110000111011011010",
		b"11111111110000111010110111",
		b"11111111110000111010110100",
		b"11111111110000111011010010",
		b"11111111110000111100010001",
		b"11111111110000111101101111",
		b"11111111110000111111101110",
		b"11111111110001000010001101",
		b"11111111110001000101001100",
		b"11111111110001001000101010",
		b"11111111110001001100101000",
		b"11111111110001010001000101",
		b"11111111110001010110000001",
		b"11111111110001011011011011",
		b"11111111110001100001010011",
		b"11111111110001100111101010",
		b"11111111110001101110011110",
		b"11111111110001110101101111",
		b"11111111110001111101011101",
		b"11111111110010000101101000",
		b"11111111110010001110001111",
		b"11111111110010010111010001",
		b"11111111110010100000101111",
		b"11111111110010101010101000",
		b"11111111110010110100111100",
		b"11111111110010111111101010",
		b"11111111110011001010110001",
		b"11111111110011010110010001",
		b"11111111110011100010001010",
		b"11111111110011101110011100",
		b"11111111110011111011000101",
		b"11111111110100001000000101",
		b"11111111110100010101011100",
		b"11111111110100100011001000",
		b"11111111110100110001001011",
		b"11111111110100111111100010",
		b"11111111110101001110001110",
		b"11111111110101011101001110",
		b"11111111110101101100100001",
		b"11111111110101111100000111",
		b"11111111110110001011111111",
		b"11111111110110011100001000",
		b"11111111110110101100100011",
		b"11111111110110111101001101",
		b"11111111110111001110001000",
		b"11111111110111011111010001",
		b"11111111110111110000101001",
		b"11111111111000000010001110",
		b"11111111111000010100000001",
		b"11111111111000100110000000",
		b"11111111111000111000001011",
		b"11111111111001001010100010",
		b"11111111111001011101000010",
		b"11111111111001101111101101",
		b"11111111111010000010100001",
		b"11111111111010010101011101",
		b"11111111111010101000100001",
		b"11111111111010111011101101",
		b"11111111111011001110111111",
		b"11111111111011100010010111",
		b"11111111111011110101110100",
		b"11111111111100001001010101",
		b"11111111111100011100111011",
		b"11111111111100110000100011",
		b"11111111111101000100001110",
		b"11111111111101010111111011",
		b"11111111111101101011101001",
		b"11111111111101111111011000",
		b"11111111111110010011000110",
		b"11111111111110100110110100",
		b"11111111111110111010100000",
		b"11111111111111001110001001",
		b"11111111111111100001110000",
		b"11111111111111110101010100",
		b"00000000000000001000110100",
		b"00000000000000011100001110",
		b"00000000000000101111100100",
		b"00000000000001000010110011",
		b"00000000000001010101111100",
		b"00000000000001101000111110",
		b"00000000000001111011110111",
		b"00000000000010001110101000",
		b"00000000000010100001010001",
		b"00000000000010110011101111",
		b"00000000000011000110000100",
		b"00000000000011011000001101",
		b"00000000000011101010001011",
		b"00000000000011111011111110",
		b"00000000000100001101100011",
		b"00000000000100011110111100",
		b"00000000000100110000000111",
		b"00000000000101000001000100",
		b"00000000000101010001110011",
		b"00000000000101100010010010",
		b"00000000000101110010100010",
		b"00000000000110000010100001",
		b"00000000000110010010010000",
		b"00000000000110100001101110",
		b"00000000000110110000111011",
		b"00000000000110111111110101",
		b"00000000000111001110011110",
		b"00000000000111011100110011",
		b"00000000000111101010110101",
		b"00000000000111111000100100",
		b"00000000001000000101111110",
		b"00000000001000010011000101",
		b"00000000001000011111110110",
		b"00000000001000101100010010",
		b"00000000001000111000011001",
		b"00000000001001000100001011",
		b"00000000001001001111100110",
		b"00000000001001011010101011",
		b"00000000001001100101011001",
		b"00000000001001101111110000",
		b"00000000001001111001110000",
		b"00000000001010000011011000",
		b"00000000001010001100101001",
		b"00000000001010010101100010",
		b"00000000001010011110000011",
		b"00000000001010100110001011",
		b"00000000001010101101111011",
		b"00000000001010110101010011",
		b"00000000001010111100010001",
		b"00000000001011000010110111",
		b"00000000001011001001000011",
		b"00000000001011001110110110",
		b"00000000001011010100010000",
		b"00000000001011011001010001",
		b"00000000001011011101110111",
		b"00000000001011100010000101",
		b"00000000001011100101111001",
		b"00000000001011101001010011",
		b"00000000001011101100010100",
		b"00000000001011101110111010",
		b"00000000001011110001001000",
		b"00000000001011110010111011",
		b"00000000001011110100010101",
		b"00000000001011110101010110",
		b"00000000001011110101111101",
		b"00000000001011110110001010",
		b"00000000001011110101111110",
		b"00000000001011110101011001",
		b"00000000001011110100011011",
		b"00000000001011110011000100",
		b"00000000001011110001010100",
		b"00000000001011101111001011",
		b"00000000001011101100101001",
		b"00000000001011101001110000",
		b"00000000001011100110011110",
		b"00000000001011100010110011",
		b"00000000001011011110110010",
		b"00000000001011011010011000",
		b"00000000001011010101100111",
		b"00000000001011010000011111",
		b"00000000001011001011000000",
		b"00000000001011000101001011",
		b"00000000001010111110111111",
		b"00000000001010111000011101",
		b"00000000001010110001100110",
		b"00000000001010101010011000",
		b"00000000001010100010110110",
		b"00000000001010011010111111",
		b"00000000001010010010110100",
		b"00000000001010001010010100",
		b"00000000001010000001100001",
		b"00000000001001111000011010",
		b"00000000001001101111000000",
		b"00000000001001100101010011",
		b"00000000001001011011010100",
		b"00000000001001010001000100",
		b"00000000001001000110100001",
		b"00000000001000111011101110",
		b"00000000001000110000101010",
		b"00000000001000100101010110",
		b"00000000001000011001110010",
		b"00000000001000001101111111",
		b"00000000001000000001111100",
		b"00000000000111110101101011",
		b"00000000000111101001001101",
		b"00000000000111011100100000",
		b"00000000000111001111100111",
		b"00000000000111000010100001",
		b"00000000000110110101001111",
		b"00000000000110100111110001",
		b"00000000000110011010001000",
		b"00000000000110001100010100",
		b"00000000000101111110010111",
		b"00000000000101110000001111",
		b"00000000000101100001111110",
		b"00000000000101010011100101",
		b"00000000000101000101000011",
		b"00000000000100110110011010",
		b"00000000000100100111101010",
		b"00000000000100011000110011",
		b"00000000000100001001110101",
		b"00000000000011111010110011",
		b"00000000000011101011101011",
		b"00000000000011011100011110",
		b"00000000000011001101001110",
		b"00000000000010111101111001",
		b"00000000000010101110100010",
		b"00000000000010011111001000",
		b"00000000000010001111101101",
		b"00000000000010000000010000",
		b"00000000000001110000110001",
		b"00000000000001100001010011",
		b"00000000000001010001110100",
		b"00000000000001000010010110",
		b"00000000000000110010111001",
		b"00000000000000100011011101",
		b"00000000000000010100000100",
		b"00000000000000000100101101",
		b"11111111111111110101011001",
		b"11111111111111100110001001",
		b"11111111111111010110111101",
		b"11111111111111000111110101",
		b"11111111111110111000110011",
		b"11111111111110101001110101",
		b"11111111111110011010111110",
		b"11111111111110001100001101",
		b"11111111111101111101100100",
		b"11111111111101101111000001",
		b"11111111111101100000100110",
		b"11111111111101010010010100",
		b"11111111111101000100001010",
		b"11111111111100110110001001",
		b"11111111111100101000010010",
		b"11111111111100011010100101",
		b"11111111111100001101000010",
		b"11111111111011111111101010",
		b"11111111111011110010011101",
		b"11111111111011100101011100",
		b"11111111111011011000100110",
		b"11111111111011001011111101",
		b"11111111111010111111100001",
		b"11111111111010110011010010",
		b"11111111111010100111010000",
		b"11111111111010011011011100",
		b"11111111111010001111110110",
		b"11111111111010000100011111",
		b"11111111111001111001010110",
		b"11111111111001101110011101",
		b"11111111111001100011110011",
		b"11111111111001011001011001",
		b"11111111111001001111001110",
		b"11111111111001000101010100",
		b"11111111111000111011101011",
		b"11111111111000110010010010",
		b"11111111111000101001001010",
		b"11111111111000100000010100",
		b"11111111111000010111101111",
		b"11111111111000001111011011",
		b"11111111111000000111011010",
		b"11111111110111111111101011",
		b"11111111110111111000001110",
		b"11111111110111110001000100",
		b"11111111110111101010001101",
		b"11111111110111100011101000",
		b"11111111110111011101010110",
		b"11111111110111010111011000",
		b"11111111110111010001101101",
		b"11111111110111001100010101",
		b"11111111110111000111010000",
		b"11111111110111000010100000",
		b"11111111110110111110000011",
		b"11111111110110111001111010",
		b"11111111110110110110000100",
		b"11111111110110110010100011",
		b"11111111110110101111010101",
		b"11111111110110101100011100",
		b"11111111110110101001110111",
		b"11111111110110100111100101",
		b"11111111110110100101101000",
		b"11111111110110100011111111",
		b"11111111110110100010101010",
		b"11111111110110100001101000",
		b"11111111110110100000111011",
		b"11111111110110100000100010",
		b"11111111110110100000011101",
		b"11111111110110100000101011",
		b"11111111110110100001001110",
		b"11111111110110100010000100",
		b"11111111110110100011001110",
		b"11111111110110100100101011",
		b"11111111110110100110011011",
		b"11111111110110101000011111",
		b"11111111110110101010110110",
		b"11111111110110101101100000",
		b"11111111110110110000011101",
		b"11111111110110110011101101",
		b"11111111110110110111001111",
		b"11111111110110111011000011",
		b"11111111110110111111001010",
		b"11111111110111000011100011",
		b"11111111110111001000001101",
		b"11111111110111001101001010",
		b"11111111110111010010010111",
		b"11111111110111010111110110",
		b"11111111110111011101100110",
		b"11111111110111100011100110",
		b"11111111110111101001110111",
		b"11111111110111110000011000",
		b"11111111110111110111001001",
		b"11111111110111111110001010",
		b"11111111111000000101011010",
		b"11111111111000001100111001",
		b"11111111111000010100100111",
		b"11111111111000011100100100",
		b"11111111111000100100101110",
		b"11111111111000101101000111",
		b"11111111111000110101101110",
		b"11111111111000111110100010",
		b"11111111111001000111100010",
		b"11111111111001010000110000",
		b"11111111111001011010001010",
		b"11111111111001100011101111",
		b"11111111111001101101100001",
		b"11111111111001110111011110",
		b"11111111111010000001100101",
		b"11111111111010001011111000",
		b"11111111111010010110010100",
		b"11111111111010100000111011",
		b"11111111111010101011101011",
		b"11111111111010110110100100",
		b"11111111111011000001100110",
		b"11111111111011001100110000",
		b"11111111111011011000000010",
		b"11111111111011100011011100",
		b"11111111111011101110111110",
		b"11111111111011111010100110",
		b"11111111111100000110010100",
		b"11111111111100010010001001",
		b"11111111111100011110000011",
		b"11111111111100101010000011",
		b"11111111111100110110000111",
		b"11111111111101000010010000",
		b"11111111111101001110011101",
		b"11111111111101011010101110",
		b"11111111111101100111000010",
		b"11111111111101110011011001",
		b"11111111111101111111110011",
		b"11111111111110001100001110",
		b"11111111111110011000101100",
		b"11111111111110100101001010",
		b"11111111111110110001101010",
		b"11111111111110111110001010",
		b"11111111111111001010101010",
		b"11111111111111010111001010",
		b"11111111111111100011101001",
		b"11111111111111110000001000",
		b"11111111111111111100100100",
		b"00000000000000001000111111",
		b"00000000000000010101011000",
		b"00000000000000100001101110",
		b"00000000000000101110000001",
		b"00000000000000111010010001",
		b"00000000000001000110011101",
		b"00000000000001010010100101",
		b"00000000000001011110101001",
		b"00000000000001101010100111",
		b"00000000000001110110100001",
		b"00000000000010000010010101",
		b"00000000000010001110000011",
		b"00000000000010011001101010",
		b"00000000000010100101001011",
		b"00000000000010110000100101",
		b"00000000000010111011111000",
		b"00000000000011000111000011",
		b"00000000000011010010000111",
		b"00000000000011011101000010",
		b"00000000000011100111110100",
		b"00000000000011110010011110",
		b"00000000000011111100111110",
		b"00000000000100000111010101",
		b"00000000000100010001100010",
		b"00000000000100011011100100",
		b"00000000000100100101011101",
		b"00000000000100101111001011",
		b"00000000000100111000101101",
		b"00000000000101000010000101",
		b"00000000000101001011010001",
		b"00000000000101010100010010",
		b"00000000000101011101000110",
		b"00000000000101100101101110",
		b"00000000000101101110001010",
		b"00000000000101110110011001",
		b"00000000000101111110011100",
		b"00000000000110000110010001",
		b"00000000000110001101111001",
		b"00000000000110010101010011",
		b"00000000000110011100011111",
		b"00000000000110100011011110",
		b"00000000000110101010001111",
		b"00000000000110110000110001",
		b"00000000000110110111000101",
		b"00000000000110111101001010",
		b"00000000000111000011000001",
		b"00000000000111001000101001",
		b"00000000000111001110000001",
		b"00000000000111010011001011",
		b"00000000000111011000000101",
		b"00000000000111011100110000",
		b"00000000000111100001001100",
		b"00000000000111100101011000",
		b"00000000000111101001010100",
		b"00000000000111101101000001",
		b"00000000000111110000011101",
		b"00000000000111110011101010",
		b"00000000000111110110100111",
		b"00000000000111111001010100",
		b"00000000000111111011110001",
		b"00000000000111111101111110",
		b"00000000000111111111111010",
		b"00000000001000000001100111",
		b"00000000001000000011000011",
		b"00000000001000000100010000",
		b"00000000001000000101001100",
		b"00000000001000000101111000",
		b"00000000001000000110010100",
		b"00000000001000000110100000",
		b"00000000001000000110011011",
		b"00000000001000000110000111",
		b"00000000001000000101100011",
		b"00000000001000000100101111",
		b"00000000001000000011101011",
		b"00000000001000000010010111",
		b"00000000001000000000110100",
		b"00000000000111111111000000",
		b"00000000000111111100111110",
		b"00000000000111111010101100",
		b"00000000000111111000001010",
		b"00000000000111110101011010",
		b"00000000000111110010011010",
		b"00000000000111101111001011",
		b"00000000000111101011101101",
		b"00000000000111101000000001",
		b"00000000000111100100000110",
		b"00000000000111011111111100",
		b"00000000000111011011100101",
		b"00000000000111010110111111",
		b"00000000000111010010001011",
		b"00000000000111001101001010",
		b"00000000000111000111111010",
		b"00000000000111000010011110",
		b"00000000000110111100110100",
		b"00000000000110110110111101",
		b"00000000000110110000111010",
		b"00000000000110101010101001",
		b"00000000000110100100001101",
		b"00000000000110011101100100",
		b"00000000000110010110101111",
		b"00000000000110001111101110",
		b"00000000000110001000100010",
		b"00000000000110000001001011",
		b"00000000000101111001101000",
		b"00000000000101110001111011",
		b"00000000000101101010000011",
		b"00000000000101100010000001",
		b"00000000000101011001110100",
		b"00000000000101010001011110",
		b"00000000000101001000111111",
		b"00000000000101000000010110",
		b"00000000000100110111100100",
		b"00000000000100101110101010",
		b"00000000000100100101100111",
		b"00000000000100011100011100",
		b"00000000000100010011001001",
		b"00000000000100001001101110",
		b"00000000000100000000001100",
		b"00000000000011110110100011",
		b"00000000000011101100110100",
		b"00000000000011100010111101",
		b"00000000000011011001000001",
		b"00000000000011001110111111",
		b"00000000000011000100111000",
		b"00000000000010111010101011",
		b"00000000000010110000011001",
		b"00000000000010100110000011",
		b"00000000000010011011101000",
		b"00000000000010010001001001",
		b"00000000000010000110100111",
		b"00000000000001111100000001",
		b"00000000000001110001011000",
		b"00000000000001100110101100",
		b"00000000000001011011111110",
		b"00000000000001010001001101",
		b"00000000000001000110011011",
		b"00000000000000111011100111",
		b"00000000000000110000110010",
		b"00000000000000100101111100",
		b"00000000000000011011000101",
		b"00000000000000010000001110",
		b"00000000000000000101010111",
		b"11111111111111111010100001",
		b"11111111111111101111101011",
		b"11111111111111100100110110",
		b"11111111111111011010000010",
		b"11111111111111001111001111",
		b"11111111111111000100011110",
		b"11111111111110111001110000",
		b"11111111111110101111000100",
		b"11111111111110100100011010",
		b"11111111111110011001110100",
		b"11111111111110001111010001",
		b"11111111111110000100110001",
		b"11111111111101111010010101",
		b"11111111111101101111111110",
		b"11111111111101100101101010",
		b"11111111111101011011011100",
		b"11111111111101010001010010",
		b"11111111111101000111001110",
		b"11111111111100111101001111",
		b"11111111111100110011010110",
		b"11111111111100101001100011",
		b"11111111111100011111110110",
		b"11111111111100010110010000",
		b"11111111111100001100110001",
		b"11111111111100000011011000",
		b"11111111111011111010000111",
		b"11111111111011110000111110",
		b"11111111111011100111111100",
		b"11111111111011011111000011",
		b"11111111111011010110010001",
		b"11111111111011001101101000",
		b"11111111111011000101001000",
		b"11111111111010111100110000",
		b"11111111111010110100100010",
		b"11111111111010101100011101",
		b"11111111111010100100100010",
		b"11111111111010011100110000",
		b"11111111111010010101001000",
		b"11111111111010001101101011",
		b"11111111111010000110010111",
		b"11111111111001111111001111",
		b"11111111111001111000010000",
		b"11111111111001110001011101",
		b"11111111111001101010110101",
		b"11111111111001100100010111",
		b"11111111111001011110000110",
		b"11111111111001010111111111",
		b"11111111111001010010000100",
		b"11111111111001001100010101",
		b"11111111111001000110110010",
		b"11111111111001000001011011",
		b"11111111111000111100010000",
		b"11111111111000110111010001",
		b"11111111111000110010011111",
		b"11111111111000101101111001",
		b"11111111111000101001011111",
		b"11111111111000100101010011",
		b"11111111111000100001010011",
		b"11111111111000011101100000",
		b"11111111111000011001111010",
		b"11111111111000010110100001",
		b"11111111111000010011010101",
		b"11111111111000010000010110",
		b"11111111111000001101100101",
		b"11111111111000001011000001",
		b"11111111111000001000101010",
		b"11111111111000000110100000",
		b"11111111111000000100100100",
		b"11111111111000000010110110",
		b"11111111111000000001010100",
		b"11111111111000000000000001",
		b"11111111110111111110111011",
		b"11111111110111111110000010",
		b"11111111110111111101010111",
		b"11111111110111111100111010",
		b"11111111110111111100101010",
		b"11111111110111111100101000",
		b"11111111110111111100110011",
		b"11111111110111111101001011",
		b"11111111110111111101110010",
		b"11111111110111111110100101",
		b"11111111110111111111100110",
		b"11111111111000000000110101",
		b"11111111111000000010010000",
		b"11111111111000000011111001",
		b"11111111111000000101110000",
		b"11111111111000000111110011",
		b"11111111111000001010000100",
		b"11111111111000001100100010",
		b"11111111111000001111001100",
		b"11111111111000010010000100",
		b"11111111111000010101001000",
		b"11111111111000011000011001",
		b"11111111111000011011110111",
		b"11111111111000011111100001",
		b"11111111111000100011011000",
		b"11111111111000100111011011",
		b"11111111111000101011101010",
		b"11111111111000110000000110",
		b"11111111111000110100101101",
		b"11111111111000111001100001",
		b"11111111111000111110100000",
		b"11111111111001000011101011",
		b"11111111111001001001000001",
		b"11111111111001001110100011",
		b"11111111111001010100010000",
		b"11111111111001011010001000",
		b"11111111111001100000001011",
		b"11111111111001100110011001",
		b"11111111111001101100110001",
		b"11111111111001110011010100",
		b"11111111111001111010000010",
		b"11111111111010000000111001",
		b"11111111111010000111111011",
		b"11111111111010001111000110",
		b"11111111111010010110011011",
		b"11111111111010011101111010",
		b"11111111111010100101100010",
		b"11111111111010101101010011",
		b"11111111111010110101001101",
		b"11111111111010111101010000",
		b"11111111111011000101011011",
		b"11111111111011001101101111",
		b"11111111111011010110001011",
		b"11111111111011011110101111",
		b"11111111111011100111011011",
		b"11111111111011110000001111",
		b"11111111111011111001001010",
		b"11111111111100000010001100",
		b"11111111111100001011010110",
		b"11111111111100010100100110",
		b"11111111111100011101111101",
		b"11111111111100100111011010",
		b"11111111111100110000111110",
		b"11111111111100111010100111",
		b"11111111111101000100010111",
		b"11111111111101001110001100",
		b"11111111111101011000000110",
		b"11111111111101100010000110",
		b"11111111111101101100001010",
		b"11111111111101110110010100",
		b"11111111111110000000100001",
		b"11111111111110001010110100",
		b"11111111111110010101001010",
		b"11111111111110011111100100",
		b"11111111111110101010000010",
		b"11111111111110110100100011",
		b"11111111111110111111001000",
		b"11111111111111001001110000",
		b"11111111111111010100011010",
		b"11111111111111011111000111",
		b"11111111111111101001110111",
		b"11111111111111110100101001",
		b"11111111111111111111011100",
		b"00000000000000001010010010",
		b"00000000000000010101001001",
		b"00000000000000100000000001",
		b"00000000000000101010111010",
		b"00000000000000110101110101",
		b"00000000000001000000110000",
		b"00000000000001001011101011",
		b"00000000000001010110100111",
		b"00000000000001100001100011",
		b"00000000000001101100011111",
		b"00000000000001110111011010",
		b"00000000000010000010010101",
		b"00000000000010001101001111",
		b"00000000000010011000001001",
		b"00000000000010100011000001",
		b"00000000000010101101110111",
		b"00000000000010111000101101",
		b"00000000000011000011100000",
		b"00000000000011001110010010",
		b"00000000000011011001000001",
		b"00000000000011100011101110",
		b"00000000000011101110011001",
		b"00000000000011111001000001",
		b"00000000000100000011100110",
		b"00000000000100001110001000",
		b"00000000000100011000100111",
		b"00000000000100100011000011",
		b"00000000000100101101011011",
		b"00000000000100110111101111",
		b"00000000000101000001111111",
		b"00000000000101001100001100",
		b"00000000000101010110010100",
		b"00000000000101100000010111",
		b"00000000000101101010010110",
		b"00000000000101110100010001",
		b"00000000000101111110000110",
		b"00000000000110000111110111",
		b"00000000000110010001100010",
		b"00000000000110011011001000",
		b"00000000000110100100101000",
		b"00000000000110101110000011",
		b"00000000000110110111011001",
		b"00000000000111000000101000",
		b"00000000000111001001110001",
		b"00000000000111010010110100",
		b"00000000000111011011110001",
		b"00000000000111100100101000",
		b"00000000000111101101011000",
		b"00000000000111110110000001",
		b"00000000000111111110100100",
		b"00000000001000000110111111",
		b"00000000001000001111010100",
		b"00000000001000010111100010",
		b"00000000001000011111101000",
		b"00000000001000100111101000",
		b"00000000001000101111011111",
		b"00000000001000110111010000",
		b"00000000001000111110111001",
		b"00000000001001000110011010",
		b"00000000001001001101110011",
		b"00000000001001010101000101",
		b"00000000001001011100001111",
		b"00000000001001100011010000",
		b"00000000001001101010001010",
		b"00000000001001110000111100",
		b"00000000001001110111100101",
		b"00000000001001111110000110",
		b"00000000001010000100011111",
		b"00000000001010001010110000",
		b"00000000001010010000111000",
		b"00000000001010010110111000",
		b"00000000001010011100101111",
		b"00000000001010100010011101",
		b"00000000001010101000000011",
		b"00000000001010101101100001",
		b"00000000001010110010110101",
		b"00000000001010111000000001",
		b"00000000001010111101000100",
		b"00000000001011000001111111",
		b"00000000001011000110110000",
		b"00000000001011001011011001",
		b"00000000001011001111111001",
		b"00000000001011010100010001",
		b"00000000001011011000011111",
		b"00000000001011011100100100",
		b"00000000001011100000100001",
		b"00000000001011100100010101",
		b"00000000001011101000000000",
		b"00000000001011101011100010",
		b"00000000001011101110111011",
		b"00000000001011110010001011",
		b"00000000001011110101010011",
		b"00000000001011111000010001",
		b"00000000001011111011000111",
		b"00000000001011111101110100",
		b"00000000001100000000011000",
		b"00000000001100000010110100",
		b"00000000001100000101000111",
		b"00000000001100000111010001",
		b"00000000001100001001010010",
		b"00000000001100001011001011",
		b"00000000001100001100111011",
		b"00000000001100001110100010",
		b"00000000001100010000000010",
		b"00000000001100010001011000",
		b"00000000001100010010100110",
		b"00000000001100010011101100",
		b"00000000001100010100101001",
		b"00000000001100010101011111",
		b"00000000001100010110001011",
		b"00000000001100010110110000",
		b"00000000001100010111001101",
		b"00000000001100010111100001",
		b"00000000001100010111101110",
		b"00000000001100010111110010",
		b"00000000001100010111101111",
		b"00000000001100010111100100",
		b"00000000001100010111010001",
		b"00000000001100010110110111",
		b"00000000001100010110010100",
		b"00000000001100010101101011",
		b"00000000001100010100111010",
		b"00000000001100010100000001",
		b"00000000001100010011000010",
		b"00000000001100010001111011",
		b"00000000001100010000101100",
		b"00000000001100001111010111",
		b"00000000001100001101111011",
		b"00000000001100001100011000",
		b"00000000001100001010101110",
		b"00000000001100001000111110",
		b"00000000001100000111000111",
		b"00000000001100000101001001",
		b"00000000001100000011000101",
		b"00000000001100000000111010",
		b"00000000001011111110101001",
		b"00000000001011111100010010",
		b"00000000001011111001110101",
		b"00000000001011110111010010",
		b"00000000001011110100101010",
		b"00000000001011110001111011",
		b"00000000001011101111000111",
		b"00000000001011101100001101",
		b"00000000001011101001001101",
		b"00000000001011100110001000",
		b"00000000001011100010111110",
		b"00000000001011011111101111",
		b"00000000001011011100011010",
		b"00000000001011011001000001",
		b"00000000001011010101100011",
		b"00000000001011010010000000",
		b"00000000001011001110011000",
		b"00000000001011001010101100",
		b"00000000001011000110111011",
		b"00000000001011000011000110",
		b"00000000001010111111001100",
		b"00000000001010111011001110",
		b"00000000001010110111001101",
		b"00000000001010110011000111",
		b"00000000001010101110111101",
		b"00000000001010101010110000",
		b"00000000001010100110011111",
		b"00000000001010100010001011",
		b"00000000001010011101110011",
		b"00000000001010011001010111",
		b"00000000001010010100111001",
		b"00000000001010010000010111",
		b"00000000001010001011110011",
		b"00000000001010000111001011",
		b"00000000001010000010100000",
		b"00000000001001111101110011",
		b"00000000001001111001000011",
		b"00000000001001110100010001",
		b"00000000001001101111011100",
		b"00000000001001101010100101",
		b"00000000001001100101101100",
		b"00000000001001100000110000",
		b"00000000001001011011110010",
		b"00000000001001010110110011",
		b"00000000001001010001110010",
		b"00000000001001001100101110",
		b"00000000001001000111101010",
		b"00000000001001000010100011",
		b"00000000001000111101011100",
		b"00000000001000111000010010",
		b"00000000001000110011001000",
		b"00000000001000101101111100",
		b"00000000001000101000110000",
		b"00000000001000100011100010",
		b"00000000001000011110010011",
		b"00000000001000011001000100",
		b"00000000001000010011110100",
		b"00000000001000001110100011",
		b"00000000001000001001010001",
		b"00000000001000000011111111",
		b"00000000000111111110101101",
		b"00000000000111111001011010",
		b"00000000000111110100000111",
		b"00000000000111101110110100",
		b"00000000000111101001100001",
		b"00000000000111100100001110",
		b"00000000000111011110111011",
		b"00000000000111011001101000",
		b"00000000000111010100010101",
		b"00000000000111001111000011",
		b"00000000000111001001110001",
		b"00000000000111000100011111",
		b"00000000000110111111001110",
		b"00000000000110111001111110",
		b"00000000000110110100101110",
		b"00000000000110101111011111",
		b"00000000000110101010010000",
		b"00000000000110100101000011",
		b"00000000000110011111110110",
		b"00000000000110011010101011",
		b"00000000000110010101100000",
		b"00000000000110010000010111",
		b"00000000000110001011001110",
		b"00000000000110000110000111",
		b"00000000000110000001000001",
		b"00000000000101111011111101",
		b"00000000000101110110111010",
		b"00000000000101110001111000",
		b"00000000000101101100111000",
		b"00000000000101100111111001",
		b"00000000000101100010111100",
		b"00000000000101011110000001",
		b"00000000000101011001000111",
		b"00000000000101010100001111",
		b"00000000000101001111011001",
		b"00000000000101001010100100",
		b"00000000000101000101110010",
		b"00000000000101000001000001",
		b"00000000000100111100010011",
		b"00000000000100110111100110",
		b"00000000000100110010111011",
		b"00000000000100101110010010",
		b"00000000000100101001101100",
		b"00000000000100100101000111",
		b"00000000000100100000100101",
		b"00000000000100011100000101",
		b"00000000000100010111100111",
		b"00000000000100010011001011",
		b"00000000000100001110110010",
		b"00000000000100001010011011",
		b"00000000000100000110000110",
		b"00000000000100000001110100",
		b"00000000000011111101100100",
		b"00000000000011111001010110",
		b"00000000000011110101001011",
		b"00000000000011110001000010",
		b"00000000000011101100111100",
		b"00000000000011101000111000",
		b"00000000000011100100110110",
		b"00000000000011100000111000",
		b"00000000000011011100111011",
		b"00000000000011011001000001",
		b"00000000000011010101001010",
		b"00000000000011010001010110",
		b"00000000000011001101100100",
		b"00000000000011001001110100",
		b"00000000000011000110000111",
		b"00000000000011000010011101",
		b"00000000000010111110110101",
		b"00000000000010111011010000",
		b"00000000000010110111101110",
		b"00000000000010110100001110",
		b"00000000000010110000110001",
		b"00000000000010101101010110",
		b"00000000000010101001111110",
		b"00000000000010100110101001",
		b"00000000000010100011010110",
		b"00000000000010100000000110",
		b"00000000000010011100111001",
		b"00000000000010011001101110",
		b"00000000000010010110100110",
		b"00000000000010010011100001",
		b"00000000000010010000011110",
		b"00000000000010001101011110",
		b"00000000000010001010100000",
		b"00000000000010000111100101",
		b"00000000000010000100101101",
		b"00000000000010000001110111",
		b"00000000000001111111000100",
		b"00000000000001111100010100",
		b"00000000000001111001100110",
		b"00000000000001110110111010",
		b"00000000000001110100010001",
		b"00000000000001110001101011",
		b"00000000000001101111000111",
		b"00000000000001101100100110",
		b"00000000000001101010000111",
		b"00000000000001100111101011",
		b"00000000000001100101010001",
		b"00000000000001100010111001",
		b"00000000000001100000100100",
		b"00000000000001011110010010",
		b"00000000000001011100000010",
		b"00000000000001011001110100",
		b"00000000000001010111101001",
		b"00000000000001010101100000",
		b"00000000000001010011011001",
		b"00000000000001010001010101",
		b"00000000000001001111010011",
		b"00000000000001001101010011",
		b"00000000000001001011010110",
		b"00000000000001001001011010",
		b"00000000000001000111100001",
		b"00000000000001000101101011",
		b"00000000000001000011110110",
		b"00000000000001000010000100",
		b"00000000000001000000010100",
		b"00000000000000111110100101",
		b"00000000000000111100111001",
		b"00000000000000111011010000",
		b"00000000000000111001101000",
		b"00000000000000111000000010",
		b"00000000000000110110011110",
		b"00000000000000110100111100",
		b"00000000000000110011011101",
		b"00000000000000110001111111",
		b"00000000000000110000100011",
		b"00000000000000101111001001",
		b"00000000000000101101110001",
		b"00000000000000101100011011",
		b"00000000000000101011000110",
		b"00000000000000101001110100",
		b"00000000000000101000100011",
		b"00000000000000100111010100",
		b"00000000000000100110000111",
		b"00000000000000100100111011",
		b"00000000000000100011110001",
		b"00000000000000100010101001",
		b"00000000000000100001100011",
		b"00000000000000100000011110",
		b"00000000000000011111011010",
		b"00000000000000011110011001",
		b"00000000000000011101011001",
		b"00000000000000011100011010",
		b"00000000000000011011011101",
		b"00000000000000011010100001",
		b"00000000000000011001100111",
		b"00000000000000011000101111",
		b"00000000000000010111110111",
		b"00000000000000010111000010",
		b"00000000000000010110001101",
		b"00000000000000010101011010",
		b"00000000000000010100101000",
		b"00000000000000010011111000",
		b"00000000000000010011001001",
		b"00000000000000010010011011",
		b"00000000000000010001101110",
		b"00000000000000010001000010",
		b"00000000000000010000011000",
		b"00000000000000001111101111",
		b"00000000000000001111000111",
		b"00000000000000001110100000",
		b"00000000000000001101111011",
		b"00000000000000001101010110",
		b"00000000000000001100110010",
		b"00000000000000001100010000",
		b"00000000000000001011101110",
		b"00000000000000001011001110",
		b"00000000000000001010101110",
		b"00000000000000001010010000",
		b"00000000000000001001110010",
		b"00000000000000001001010110",
		b"00000000000000001000111010",
		b"00000000000000001000011111",
		b"00000000000000001000000101",
		b"00000000000000000111101100",
		b"00000000000000000111010100",
		b"00000000000000000110111100",
		b"00000000000000000110100101",
		b"00000000000000000110001111",
		b"00000000000000000101111010",
		b"00000000000000000101100110",
		b"00000000000000000101010010",
		b"00000000000000000100111111",
		b"00000000000000000100101100",
		b"00000000000000000100011011",
		b"00000000000000000100001010",
		b"00000000000000000011111001",
		b"00000000000000000011101010",
		b"00000000000000000011011010",
		b"00000000000000000011001100",
		b"00000000000000000010111110",
		b"00000000000000000010110000",
		b"00000000000000000010100011",
		b"00000000000000000010010111",
		b"00000000000000000010001011",
		b"00000000000000000010000000",
		b"00000000000000000001110101",
		b"00000000000000000001101010",
		b"00000000000000000001100000",
		b"00000000000000000001010111",
		b"00000000000000000001001110",
		b"00000000000000000001000101",
		b"00000000000000000000111101",
		b"00000000000000000000110101",
		b"00000000000000000000101110",
		b"00000000000000000000100110",
		b"00000000000000000000100000",
		b"00000000000000000000011001",
		b"00000000000000000000010011",
		b"00000000000000000000001110",
		b"00000000000000000000001000",
		b"00000000000000000000000011",
		b"11111111111111111111111110",
		b"11111111111111111111111010",
		b"11111111111111111111110101",
		b"11111111111111111111110001",
		b"11111111111111111111101101",
		b"11111111111111111111101010",
		b"11111111111111111111100111",
		b"11111111111111111111100100",
		b"11111111111111111111100001",
		b"11111111111111111111011110",
		b"11111111111111111111011100",
		b"11111111111111111111011010",
		b"11111111111111111111010111",
		b"11111111111111111111010110",
		b"11111111111111111111010100",
		b"11111111111111111111010010",
		b"11111111111111111111010001",
		b"11111111111111111111010000",
		b"11111111111111111111001111",
		b"11111111111111111111001110",
		b"11111111111111111111001101",
		b"11111111111111111111001100",
		b"11111111111111111111001100",
		b"11111111111111111111001011",
		b"11111111111111111111001011",
		b"11111111111111111111001011",
		b"11111111111111111111001010",
		b"11111111111111111111001010",
		b"11111111111111111111001010",
		b"11111111111111111111001010",
		b"11111111111111111111001011",
		b"11111111111111111111001011",
		b"11111111111111111111001011",
		b"11111111111111111111001100",
		b"11111111111111111111001100",
		b"11111111111111111111001101",
		b"11111111111111111111001101",
		b"11111111111111111111001110",
		b"11111111111111111111001110",
		b"11111111111111111111001111",
		b"11111111111111111111010000",
		b"11111111111111111111010000",
		b"11111111111111111111010001",
		b"11111111111111111111010010",
		b"11111111111111111111010011",
		b"11111111111111111111010100",
		b"11111111111111111111010101",
		b"11111111111111111111010110",
		b"11111111111111111111010110",
		b"11111111111111111111010111",
		b"11111111111111111111011000",
		b"11111111111111111111011001",
		b"11111111111111111111011010",
		b"11111111111111111111011011",
		b"11111111111111111111011100",
		b"11111111111111111111011101",
		b"11111111111111111111011110",
		b"11111111111111111111011111",
		b"11111111111111111111100000",
		b"11111111111111111111100001",
		b"11111111111111111111100010",
		b"11111111111111111111100011",
		b"11111111111111111111100100",
		b"11111111111111111111100101",
		b"11111111111111111111100110",
		b"11111111111111111111100111",
		b"11111111111111111111101000",
		b"11111111111111111111101000",
		b"11111111111111111111101001",
		b"11111111111111111111101010",
		b"11111111111111111111101011",
		b"11111111111111111111101100",
		b"11111111111111111111101100",
		b"11111111111111111111101101",
		b"11111111111111111111101110",
		b"11111111111111111111101111",
		b"11111111111111111111101111",
		b"11111111111111111111110000",
		b"11111111111111111111110001",
		b"11111111111111111111110001",
		b"11111111111111111111110010",
		b"11111111111111111111110011",
		b"11111111111111111111110011",
		b"11111111111111111111110100",
		b"11111111111111111111110101",
		b"11111111111111111111110101",
		b"11111111111111111111110110",
		b"11111111111111111111110110",
		b"11111111111111111111110111",
		b"11111111111111111111111000",
		b"11111111111111111111111000",
		b"11111111111111111111111001",
		b"11111111111111111111111001",
		b"11111111111111111111111010",
		b"11111111111111111111111011",
		b"11111111111111111111111011",
		b"11111111111111111111111100",
		b"11111111111111111111111100",
		b"11111111111111111111111101",
		b"11111111111111111111111101",
		b"11111111111111111111111110",
		b"11111111111111111111111110",
		b"11111111111111111111111110",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000"
	);

end src_rom_pkg;