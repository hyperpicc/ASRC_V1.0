library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package src_rom_pkg is

	constant COE_WIDTH	: integer := 22;
	constant COE_CENTRE	: signed( 21 downto 0 ) := b"0111111101011100001010";

	type COE_ROM_TYPE is array( 4095 downto 0 ) of signed( 21 downto 0 );
	constant COE_ROM	 : COE_ROM_TYPE := (
		b"0111111101011001000110",
		b"0111111101001111111001",
		b"0111111101000000100100",
		b"0111111100101011000111",
		b"0111111100001111100011",
		b"0111111011101101110111",
		b"0111111011000110000110",
		b"0111111010011000001111",
		b"0111111001100100010100",
		b"0111111000101010010101",
		b"0111110111101010010101",
		b"0111110110100100010100",
		b"0111110101011000010101",
		b"0111110100000110011000",
		b"0111110010101110011111",
		b"0111110001010000101101",
		b"0111101111101101000011",
		b"0111101110000011100011",
		b"0111101100010100010001",
		b"0111101010011111001101",
		b"0111101000100100011100",
		b"0111100110100011111111",
		b"0111100100011101111001",
		b"0111100010010010001101",
		b"0111100000000000111110",
		b"0111011101101010001111",
		b"0111011011001110000100",
		b"0111011000101100100000",
		b"0111010110000101100110",
		b"0111010011011001011010",
		b"0111010000101000000000",
		b"0111001101110001011011",
		b"0111001010110101110000",
		b"0111000111110101000010",
		b"0111000100101111010110",
		b"0111000001100100101111",
		b"0110111110010101010011",
		b"0110111011000001000101",
		b"0110110111101000001011",
		b"0110110100001010101000",
		b"0110110000101000100001",
		b"0110101101000001111100",
		b"0110101001010110111110",
		b"0110100101100111101010",
		b"0110100001110100000111",
		b"0110011101111100011001",
		b"0110011010000000100110",
		b"0110010110000000110011",
		b"0110010001111101000110",
		b"0110001101110101100100",
		b"0110001001101010010010",
		b"0110000101011011010110",
		b"0110000001001000110111",
		b"0101111100110010111001",
		b"0101111000011001100010",
		b"0101110011111100111001",
		b"0101101111011101000100",
		b"0101101010111010001000",
		b"0101100110010100001011",
		b"0101100001101011010100",
		b"0101011100111111101001",
		b"0101011000010001001111",
		b"0101010011100000001110",
		b"0101001110101100101100",
		b"0101001001110110101111",
		b"0101000100111110011100",
		b"0101000000000011111100",
		b"0100111011000111010100",
		b"0100110110001000101011",
		b"0100110001001000000111",
		b"0100101100000101101111",
		b"0100100111000001101001",
		b"0100100001111011111100",
		b"0100011100110100101111",
		b"0100010111101100001000",
		b"0100010010100010001110",
		b"0100001101010111000111",
		b"0100001000001010111011",
		b"0100000010111101101111",
		b"0011111101101111101011",
		b"0011111000100000110101",
		b"0011110011010001010100",
		b"0011101110000001001110",
		b"0011101000110000101010",
		b"0011100011011111101111",
		b"0011011110001110100100",
		b"0011011000111101001110",
		b"0011010011101011110101",
		b"0011001110011010011111",
		b"0011001001001001010011",
		b"0011000011111000010111",
		b"0010111110100111110010",
		b"0010111001010111101010",
		b"0010110100001000000101",
		b"0010101110111001001010",
		b"0010101001101011000000",
		b"0010100100011101101101",
		b"0010011111010001010110",
		b"0010011010000110000010",
		b"0010010100111011111000",
		b"0010001111110010111101",
		b"0010001010101011011000",
		b"0010000101100101001110",
		b"0010000000100000100110",
		b"0001111011011101100110",
		b"0001110110011100010011",
		b"0001110001011100110010",
		b"0001101100011111001011",
		b"0001100111100011100010",
		b"0001100010101001111101",
		b"0001011101110010100010",
		b"0001011000111101010110",
		b"0001010100001010011111",
		b"0001001111011010000001",
		b"0001001010101100000010",
		b"0001000110000000100111",
		b"0001000001010111110101",
		b"0000111100110001110001",
		b"0000111000001110100001",
		b"0000110011101110001000",
		b"0000101111010000101011",
		b"0000101010110110010000",
		b"0000100110011110111010",
		b"0000100010001010101111",
		b"0000011101111001110010",
		b"0000011001101100001000",
		b"0000010101100001110100",
		b"0000010001011010111011",
		b"0000001101010111100010",
		b"0000001001010111101011",
		b"0000000101011011011010",
		b"0000000001100010110100",
		b"1111111101101101111011",
		b"1111111001111100110011",
		b"1111110110001111011111",
		b"1111110010100110000011",
		b"1111101111000000100010",
		b"1111101011011110111110",
		b"1111101000000001011011",
		b"1111100100100111111100",
		b"1111100001010010100010",
		b"1111011110000001010001",
		b"1111011010110100001011",
		b"1111010111101011010011",
		b"1111010100100110101010",
		b"1111010001100110010010",
		b"1111001110101010001110",
		b"1111001011110010100000",
		b"1111001000111111001001",
		b"1111000110010000001011",
		b"1111000011100101101000",
		b"1111000000111111100000",
		b"1110111110011101110101",
		b"1110111100000000101001",
		b"1110111001100111111100",
		b"1110110111010011101111",
		b"1110110101000100000100",
		b"1110110010111000111010",
		b"1110110000110010010010",
		b"1110101110110000001110",
		b"1110101100110010101101",
		b"1110101010111001101111",
		b"1110101001000101010101",
		b"1110100111010101011110",
		b"1110100101101010001011",
		b"1110100100000011011011",
		b"1110100010100001001110",
		b"1110100001000011100100",
		b"1110011111101010011100",
		b"1110011110010101110101",
		b"1110011101000101101111",
		b"1110011011111010001000",
		b"1110011010110011000000",
		b"1110011001110000010110",
		b"1110011000110010001000",
		b"1110010111111000010101",
		b"1110010111000010111100",
		b"1110010110010001111011",
		b"1110010101100101010000",
		b"1110010100111100111011",
		b"1110010100011000111000",
		b"1110010011111001000110",
		b"1110010011011101100100",
		b"1110010011000110001110",
		b"1110010010110011000011",
		b"1110010010100100000001",
		b"1110010010011001000101",
		b"1110010010010010001100",
		b"1110010010001111010100",
		b"1110010010010000011010",
		b"1110010010010101011101",
		b"1110010010011110010111",
		b"1110010010101011001000",
		b"1110010010111011101011",
		b"1110010011001111111110",
		b"1110010011100111111110",
		b"1110010100000011100111",
		b"1110010100100010110110",
		b"1110010101000101101000",
		b"1110010101101011111001",
		b"1110010110010101100101",
		b"1110010111000010101010",
		b"1110010111110011000011",
		b"1110011000100110101101",
		b"1110011001011101100100",
		b"1110011010010111100100",
		b"1110011011010100101001",
		b"1110011100010100101111",
		b"1110011101010111110011",
		b"1110011110011101101111",
		b"1110011111100110100001",
		b"1110100000110010000100",
		b"1110100010000000010011",
		b"1110100011010001001011",
		b"1110100100100100100111",
		b"1110100101111010100011",
		b"1110100111010010111011",
		b"1110101000101101101001",
		b"1110101010001010101010",
		b"1110101011101001111001",
		b"1110101101001011010010",
		b"1110101110101110110000",
		b"1110110000010100001111",
		b"1110110001111011101010",
		b"1110110011100100111100",
		b"1110110101010000000001",
		b"1110110110111100110100",
		b"1110111000101011010001",
		b"1110111010011011010011",
		b"1110111100001100110101",
		b"1110111101111111110010",
		b"1110111111110100000111",
		b"1111000001101001101101",
		b"1111000011100000100010",
		b"1111000101011000011111",
		b"1111000111010001100000",
		b"1111001001001011100001",
		b"1111001011000110011101",
		b"1111001101000010001111",
		b"1111001110111110110011",
		b"1111010000111100000011",
		b"1111010010111001111100",
		b"1111010100111000011000",
		b"1111010110110111010100",
		b"1111011000110110101010",
		b"1111011010110110010111",
		b"1111011100110110010100",
		b"1111011110110110011111",
		b"1111100000110110110011",
		b"1111100010110111001010",
		b"1111100100110111100001",
		b"1111100110110111110100",
		b"1111101000110111111110",
		b"1111101010110111111010",
		b"1111101100110111100110",
		b"1111101110110110111011",
		b"1111110000110101110111",
		b"1111110010110100010100",
		b"1111110100110010010000",
		b"1111110110101111100101",
		b"1111111000101100010001",
		b"1111111010101000001110",
		b"1111111100100011011010",
		b"1111111110011101110000",
		b"0000000000010111001101",
		b"0000000010001111101100",
		b"0000000100000111001011",
		b"0000000101111101100101",
		b"0000000111110010111000",
		b"0000001001100110111111",
		b"0000001011011001110111",
		b"0000001101001011011101",
		b"0000001110111011101110",
		b"0000010000101010100110",
		b"0000010010011000000011",
		b"0000010100000100000001",
		b"0000010101101110011101",
		b"0000010111010111010100",
		b"0000011000111110100100",
		b"0000011010100100001001",
		b"0000011100001000000001",
		b"0000011101101010001010",
		b"0000011111001010100000",
		b"0000100000101001000001",
		b"0000100010000101101100",
		b"0000100011100000011101",
		b"0000100100111001010010",
		b"0000100110010000001001",
		b"0000100111100101000000",
		b"0000101000110111110110",
		b"0000101010001000100111",
		b"0000101011010111010010",
		b"0000101100100011110111",
		b"0000101101101110010001",
		b"0000101110110110100001",
		b"0000101111111100100101",
		b"0000110001000000011011",
		b"0000110010000010000001",
		b"0000110011000001011000",
		b"0000110011111110011100",
		b"0000110100111001001110",
		b"0000110101110001101101",
		b"0000110110100111110110",
		b"0000110111011011101010",
		b"0000111000001101001000",
		b"0000111000111100001111",
		b"0000111001101000111110",
		b"0000111010010011010101",
		b"0000111010111011010100",
		b"0000111011100000111001",
		b"0000111100000100000110",
		b"0000111100100100111001",
		b"0000111101000011010010",
		b"0000111101011111010010",
		b"0000111101111000111001",
		b"0000111110010000000110",
		b"0000111110100100111010",
		b"0000111110110111010101",
		b"0000111111000111011000",
		b"0000111111010101000010",
		b"0000111111100000010101",
		b"0000111111101001010001",
		b"0000111111101111110111",
		b"0000111111110100001000",
		b"0000111111110110000011",
		b"0000111111110101101011",
		b"0000111111110011000000",
		b"0000111111101110000011",
		b"0000111111100110110101",
		b"0000111111011101011000",
		b"0000111111010001101100",
		b"0000111111000011110100",
		b"0000111110110011110000",
		b"0000111110100001100001",
		b"0000111110001101001010",
		b"0000111101110110101100",
		b"0000111101011110001001",
		b"0000111101000011100001",
		b"0000111100100110111000",
		b"0000111100001000001110",
		b"0000111011100111100110",
		b"0000111011000101000010",
		b"0000111010100000100011",
		b"0000111001111010001011",
		b"0000111001010001111110",
		b"0000111000100111111100",
		b"0000110111111100001000",
		b"0000110111001110100100",
		b"0000110110011111010010",
		b"0000110101101110010101",
		b"0000110100111011110000",
		b"0000110100000111100100",
		b"0000110011010001110011",
		b"0000110010011010100010",
		b"0000110001100001110001",
		b"0000110000100111100100",
		b"0000101111101011111101",
		b"0000101110101110111110",
		b"0000101101110000101011",
		b"0000101100110001000110",
		b"0000101011110000010010",
		b"0000101010101110010001",
		b"0000101001101011000110",
		b"0000101000100110110101",
		b"0000100111100001011111",
		b"0000100110011011001001",
		b"0000100101010011110011",
		b"0000100100001011100010",
		b"0000100011000010011001",
		b"0000100001111000011001",
		b"0000100000101101100111",
		b"0000011111100010000100",
		b"0000011110010101110101",
		b"0000011101001000111011",
		b"0000011011111011011010",
		b"0000011010101101010101",
		b"0000011001011110101111",
		b"0000011000001111101010",
		b"0000010111000000001010",
		b"0000010101110000010010",
		b"0000010100100000000100",
		b"0000010011001111100011",
		b"0000010001111110110011",
		b"0000010000101101110110",
		b"0000001111011100110000",
		b"0000001110001011100010",
		b"0000001100111010010001",
		b"0000001011101000111110",
		b"0000001010010111101101",
		b"0000001001000110100001",
		b"0000000111110101011100",
		b"0000000110100100100010",
		b"0000000101010011110101",
		b"0000000100000011010111",
		b"0000000010110011001100",
		b"0000000001100011010111",
		b"0000000000010011111001",
		b"1111111111000100110110",
		b"1111111101110110010001",
		b"1111111100101000001011",
		b"1111111011011010101000",
		b"1111111010001101101010",
		b"1111111001000001010100",
		b"1111110111110101101000",
		b"1111110110101010101000",
		b"1111110101100000010111",
		b"1111110100010110111000",
		b"1111110011001110001100",
		b"1111110010000110010110",
		b"1111110000111111011000",
		b"1111101111111001010101",
		b"1111101110110100001110",
		b"1111101101110000000110",
		b"1111101100101100111110",
		b"1111101011101010111010",
		b"1111101010101001111010",
		b"1111101001101010000001",
		b"1111101000101011010000",
		b"1111100111101101101010",
		b"1111100110110001010000",
		b"1111100101110110000101",
		b"1111100100111100001000",
		b"1111100100000011011110",
		b"1111100011001100000110",
		b"1111100010010110000010",
		b"1111100001100001010101",
		b"1111100000101101111110",
		b"1111011111111100000001",
		b"1111011111001011011110",
		b"1111011110011100010101",
		b"1111011101101110101010",
		b"1111011101000010011100",
		b"1111011100010111101100",
		b"1111011011101110011101",
		b"1111011011000110101110",
		b"1111011010100000100001",
		b"1111011001111011110111",
		b"1111011001011000110000",
		b"1111011000110111001101",
		b"1111011000010111001110",
		b"1111010111111000110110",
		b"1111010111011100000011",
		b"1111010111000000110111",
		b"1111010110100111010010",
		b"1111010110001111010100",
		b"1111010101111000111110",
		b"1111010101100100001111",
		b"1111010101010001001010",
		b"1111010100111111101100",
		b"1111010100101111110111",
		b"1111010100100001101011",
		b"1111010100010101000111",
		b"1111010100001010001100",
		b"1111010100000000111001",
		b"1111010011111001001110",
		b"1111010011110011001011",
		b"1111010011101110110000",
		b"1111010011101011111100",
		b"1111010011101010110000",
		b"1111010011101011001010",
		b"1111010011101101001001",
		b"1111010011110000101111",
		b"1111010011110101111001",
		b"1111010011111100100111",
		b"1111010100000100111001",
		b"1111010100001110101101",
		b"1111010100011010000100",
		b"1111010100100110111011",
		b"1111010100110101010011",
		b"1111010101000101001001",
		b"1111010101010110011110",
		b"1111010101101001010000",
		b"1111010101111101011110",
		b"1111010110010011000111",
		b"1111010110101010001001",
		b"1111010111000010100100",
		b"1111010111011100010110",
		b"1111010111110111011110",
		b"1111011000010011111010",
		b"1111011000110001101001",
		b"1111011001010000101010",
		b"1111011001110000111011",
		b"1111011010010010011011",
		b"1111011010110101001000",
		b"1111011011011001000000",
		b"1111011011111110000010",
		b"1111011100100100001101",
		b"1111011101001011011110",
		b"1111011101110011110100",
		b"1111011110011101001101",
		b"1111011111000111100111",
		b"1111011111110011000001",
		b"1111100000011111011000",
		b"1111100001001100101011",
		b"1111100001111010111001",
		b"1111100010101001111110",
		b"1111100011011001111001",
		b"1111100100001010101001",
		b"1111100100111100001010",
		b"1111100101101110011100",
		b"1111100110100001011100",
		b"1111100111010101001001",
		b"1111101000001001011111",
		b"1111101000111110011110",
		b"1111101001110100000011",
		b"1111101010101010001011",
		b"1111101011100000110110",
		b"1111101100011000000000",
		b"1111101101001111101000",
		b"1111101110000111101100",
		b"1111101111000000001001",
		b"1111101111111000111110",
		b"1111110000110010000111",
		b"1111110001101011100100",
		b"1111110010100101010010",
		b"1111110011011111001111",
		b"1111110100011001011000",
		b"1111110101010011101100",
		b"1111110110001110001001",
		b"1111110111001000101100",
		b"1111111000000011010011",
		b"1111111000111101111100",
		b"1111111001111000100101",
		b"1111111010110011001101",
		b"1111111011101101110000",
		b"1111111100101000001101",
		b"1111111101100010100001",
		b"1111111110011100101100",
		b"1111111111010110101010",
		b"0000000000010000011010",
		b"0000000001001001111001",
		b"0000000010000011000111",
		b"0000000010111100000000",
		b"0000000011110100100011",
		b"0000000100101100101101",
		b"0000000101100100011110",
		b"0000000110011011110011",
		b"0000000111010010101010",
		b"0000001000001001000001",
		b"0000001000111110111000",
		b"0000001001110100001011",
		b"0000001010101000111001",
		b"0000001011011101000000",
		b"0000001100010000100000",
		b"0000001101000011010101",
		b"0000001101110101011110",
		b"0000001110100110111011",
		b"0000001111010111101000",
		b"0000010000000111100101",
		b"0000010000110110110001",
		b"0000010001100101001001",
		b"0000010010010010101100",
		b"0000010010111111011001",
		b"0000010011101011001111",
		b"0000010100010110001100",
		b"0000010101000000001110",
		b"0000010101101001010101",
		b"0000010110010001100000",
		b"0000010110111000101101",
		b"0000010111011110111010",
		b"0000011000000100001000",
		b"0000011000101000010100",
		b"0000011001001011011111",
		b"0000011001101101100110",
		b"0000011010001110101001",
		b"0000011010101110100111",
		b"0000011011001101011111",
		b"0000011011101011010000",
		b"0000011100000111111010",
		b"0000011100100011011100",
		b"0000011100111101110101",
		b"0000011101010111000100",
		b"0000011101101111001010",
		b"0000011110000110000100",
		b"0000011110011011110100",
		b"0000011110110000010111",
		b"0000011111000011101111",
		b"0000011111010101111010",
		b"0000011111100110111000",
		b"0000011111110110101001",
		b"0000100000000101001101",
		b"0000100000010010100011",
		b"0000100000011110101011",
		b"0000100000101001100110",
		b"0000100000110011010010",
		b"0000100000111011110000",
		b"0000100001000011000001",
		b"0000100001001001000011",
		b"0000100001001101111000",
		b"0000100001010001011111",
		b"0000100001010011111000",
		b"0000100001010101000100",
		b"0000100001010101000010",
		b"0000100001010011110100",
		b"0000100001010001011010",
		b"0000100001001101110011",
		b"0000100001001001000001",
		b"0000100001000011000100",
		b"0000100000111011111100",
		b"0000100000110011101010",
		b"0000100000101010001110",
		b"0000100000011111101010",
		b"0000100000010011111101",
		b"0000100000000111001001",
		b"0000011111111001001110",
		b"0000011111101010001101",
		b"0000011111011010000110",
		b"0000011111001000111100",
		b"0000011110110110101101",
		b"0000011110100011011101",
		b"0000011110001111001010",
		b"0000011101111001110111",
		b"0000011101100011100100",
		b"0000011101001100010010",
		b"0000011100110100000011",
		b"0000011100011010111000",
		b"0000011100000000110001",
		b"0000011011100101110000",
		b"0000011011001001110110",
		b"0000011010101101000100",
		b"0000011010001111011100",
		b"0000011001110000111110",
		b"0000011001010001101100",
		b"0000011000110001101000",
		b"0000011000010000110010",
		b"0000010111101111001101",
		b"0000010111001100111001",
		b"0000010110101001110111",
		b"0000010110000110001010",
		b"0000010101100001110011",
		b"0000010100111100110010",
		b"0000010100010111001011",
		b"0000010011110000111101",
		b"0000010011001010001011",
		b"0000010010100010110110",
		b"0000010001111011000000",
		b"0000010001010010101010",
		b"0000010000101001110110",
		b"0000010000000000100101",
		b"0000001111010110111001",
		b"0000001110101100110011",
		b"0000001110000010010110",
		b"0000001101010111100011",
		b"0000001100101100011010",
		b"0000001100000000111111",
		b"0000001011010101010010",
		b"0000001010101001010110",
		b"0000001001111101001011",
		b"0000001001010000110100",
		b"0000001000100100010010",
		b"0000000111110111100110",
		b"0000000111001010110011",
		b"0000000110011101111010",
		b"0000000101110000111101",
		b"0000000101000011111100",
		b"0000000100010110111011",
		b"0000000011101001111010",
		b"0000000010111100111011",
		b"0000000010010000000000",
		b"0000000001100011001010",
		b"0000000000110110011011",
		b"0000000000001001110101",
		b"1111111111011101011000",
		b"1111111110110001000111",
		b"1111111110000101000011",
		b"1111111101011001001110",
		b"1111111100101101101001",
		b"1111111100000010010101",
		b"1111111011010111010101",
		b"1111111010101100101001",
		b"1111111010000010010011",
		b"1111111001011000010101",
		b"1111111000101110110000",
		b"1111111000000101100101",
		b"1111110111011100110101",
		b"1111110110110100100011",
		b"1111110110001100101111",
		b"1111110101100101011010",
		b"1111110100111110100111",
		b"1111110100011000010110",
		b"1111110011110010101000",
		b"1111110011001101011111",
		b"1111110010101000111100",
		b"1111110010000101000000",
		b"1111110001100001101100",
		b"1111110000111111000010",
		b"1111110000011101000010",
		b"1111101111111011101101",
		b"1111101111011011000101",
		b"1111101110111011001011",
		b"1111101110011011111111",
		b"1111101101111101100011",
		b"1111101101011111110111",
		b"1111101101000010111100",
		b"1111101100100110110100",
		b"1111101100001011011110",
		b"1111101011110000111101",
		b"1111101011010111010000",
		b"1111101010111110011000",
		b"1111101010100110010110",
		b"1111101010001111001011",
		b"1111101001111000110111",
		b"1111101001100011011011",
		b"1111101001001110111000",
		b"1111101000111011001101",
		b"1111101000101000011100",
		b"1111101000010110100101",
		b"1111101000000101101001",
		b"1111100111110101100111",
		b"1111100111100110100001",
		b"1111100111011000010110",
		b"1111100111001011000111",
		b"1111100110111110110100",
		b"1111100110110011011101",
		b"1111100110101001000011",
		b"1111100110011111100101",
		b"1111100110010111000101",
		b"1111100110001111100001",
		b"1111100110001000111010",
		b"1111100110000011010001",
		b"1111100101111110100100",
		b"1111100101111010110100",
		b"1111100101111000000010",
		b"1111100101110110001011",
		b"1111100101110101010010",
		b"1111100101110101010101",
		b"1111100101110110010100",
		b"1111100101111000010000",
		b"1111100101111011000111",
		b"1111100101111110111001",
		b"1111100110000011100110",
		b"1111100110001001001111",
		b"1111100110001111110001",
		b"1111100110010111001110",
		b"1111100110011111100011",
		b"1111100110101000110010",
		b"1111100110110010111001",
		b"1111100110111101111000",
		b"1111100111001001101110",
		b"1111100111010110011011",
		b"1111100111100011111110",
		b"1111100111110010010111",
		b"1111101000000001100011",
		b"1111101000010001100100",
		b"1111101000100010011000",
		b"1111101000110011111111",
		b"1111101001000110010111",
		b"1111101001011001011111",
		b"1111101001101101011000",
		b"1111101010000010000000",
		b"1111101010010111010110",
		b"1111101010101101011001",
		b"1111101011000100001000",
		b"1111101011011011100011",
		b"1111101011110011101000",
		b"1111101100001100010111",
		b"1111101100100101101101",
		b"1111101100111111101011",
		b"1111101101011010010000",
		b"1111101101110101011001",
		b"1111101110010001000110",
		b"1111101110101101010111",
		b"1111101111001010001001",
		b"1111101111100111011100",
		b"1111110000000101001110",
		b"1111110000100011011111",
		b"1111110001000010001100",
		b"1111110001100001010110",
		b"1111110010000000111011",
		b"1111110010100000111001",
		b"1111110011000001001111",
		b"1111110011100001111100",
		b"1111110100000010111111",
		b"1111110100100100010111",
		b"1111110101000110000010",
		b"1111110101100111111111",
		b"1111110110001010001101",
		b"1111110110101100101010",
		b"1111110111001111010101",
		b"1111110111110010001101",
		b"1111111000010101010001",
		b"1111111000111000011111",
		b"1111111001011011110110",
		b"1111111001111111010101",
		b"1111111010100010111010",
		b"1111111011000110100100",
		b"1111111011101010010010",
		b"1111111100001110000011",
		b"1111111100110001110101",
		b"1111111101010101100111",
		b"1111111101111001010111",
		b"1111111110011101000101",
		b"1111111111000000101111",
		b"1111111111100100010100",
		b"0000000000000111110010",
		b"0000000000101011001001",
		b"0000000001001110010111",
		b"0000000001110001011011",
		b"0000000010010100010011",
		b"0000000010110110111111",
		b"0000000011011001011101",
		b"0000000011111011101101",
		b"0000000100011101101100",
		b"0000000100111111011001",
		b"0000000101100000110100",
		b"0000000110000001111100",
		b"0000000110100010101111",
		b"0000000111000011001100",
		b"0000000111100011010010",
		b"0000001000000011000001",
		b"0000001000100010010110",
		b"0000001001000001010001",
		b"0000001001011111110001",
		b"0000001001111101110101",
		b"0000001010011011011100",
		b"0000001010111000100100",
		b"0000001011010101001110",
		b"0000001011110001011000",
		b"0000001100001101000000",
		b"0000001100101000001000",
		b"0000001101000010101100",
		b"0000001101011100101101",
		b"0000001101110110001010",
		b"0000001110001111000010",
		b"0000001110100111010100",
		b"0000001110111110111111",
		b"0000001111010110000011",
		b"0000001111101100011111",
		b"0000010000000010010010",
		b"0000010000010111011100",
		b"0000010000101011111100",
		b"0000010000111111110010",
		b"0000010001010010111100",
		b"0000010001100101011011",
		b"0000010001110111001101",
		b"0000010010001000010011",
		b"0000010010011000101011",
		b"0000010010101000010110",
		b"0000010010110111010011",
		b"0000010011000101100001",
		b"0000010011010011000001",
		b"0000010011011111110001",
		b"0000010011101011110010",
		b"0000010011110111000100",
		b"0000010100000001100101",
		b"0000010100001011010110",
		b"0000010100010100010111",
		b"0000010100011100100111",
		b"0000010100100100000111",
		b"0000010100101010110101",
		b"0000010100110000110011",
		b"0000010100110110000000",
		b"0000010100111010011011",
		b"0000010100111110000110",
		b"0000010101000001000000",
		b"0000010101000011001001",
		b"0000010101000100100001",
		b"0000010101000101001000",
		b"0000010101000100111110",
		b"0000010101000100000100",
		b"0000010101000010011010",
		b"0000010101000000000000",
		b"0000010100111100110110",
		b"0000010100111000111100",
		b"0000010100110100010011",
		b"0000010100101110111011",
		b"0000010100101000110101",
		b"0000010100100010000000",
		b"0000010100011010011101",
		b"0000010100010010001101",
		b"0000010100001001001111",
		b"0000010011111111100110",
		b"0000010011110101010000",
		b"0000010011101010001110",
		b"0000010011011110100010",
		b"0000010011010010001010",
		b"0000010011000101001001",
		b"0000010010110111011111",
		b"0000010010101001001100",
		b"0000010010011010010001",
		b"0000010010001010101111",
		b"0000010001111010100101",
		b"0000010001101001110110",
		b"0000010001011000100010",
		b"0000010001000110101000",
		b"0000010000110100001011",
		b"0000010000100001001011",
		b"0000010000001101101001",
		b"0000001111111001100101",
		b"0000001111100101000001",
		b"0000001111001111111101",
		b"0000001110111010011010",
		b"0000001110100100011000",
		b"0000001110001101111010",
		b"0000001101110110111111",
		b"0000001101011111101001",
		b"0000001101000111111001",
		b"0000001100101111101111",
		b"0000001100010111001100",
		b"0000001011111110010001",
		b"0000001011100101000000",
		b"0000001011001011011010",
		b"0000001010110001011110",
		b"0000001010010111001111",
		b"0000001001111100101101",
		b"0000001001100001111010",
		b"0000001001000110110101",
		b"0000001000101011100001",
		b"0000001000001111111111",
		b"0000000111110100001111",
		b"0000000111011000010010",
		b"0000000110111100001001",
		b"0000000110011111110111",
		b"0000000110000011011010",
		b"0000000101100110110110",
		b"0000000101001010001010",
		b"0000000100101101010111",
		b"0000000100010000100000",
		b"0000000011110011100100",
		b"0000000011010110100101",
		b"0000000010111001100100",
		b"0000000010011100100010",
		b"0000000001111111100000",
		b"0000000001100010011111",
		b"0000000001000101100000",
		b"0000000000101000100100",
		b"0000000000001011101100",
		b"1111111111101110111001",
		b"1111111111010010001101",
		b"1111111110110101100111",
		b"1111111110011001001010",
		b"1111111101111100110110",
		b"1111111101100000101101",
		b"1111111101000100101110",
		b"1111111100101000111100",
		b"1111111100001101010110",
		b"1111111011110001111111",
		b"1111111011010110110110",
		b"1111111010111011111110",
		b"1111111010100001010110",
		b"1111111010000111000000",
		b"1111111001101100111100",
		b"1111111001010011001100",
		b"1111111000111001110001",
		b"1111111000100000101010",
		b"1111111000000111111010",
		b"1111110111101111100000",
		b"1111110111010111011110",
		b"1111110110111111110101",
		b"1111110110101000100101",
		b"1111110110010001101110",
		b"1111110101111011010011",
		b"1111110101100101010011",
		b"1111110101001111101111",
		b"1111110100111010101000",
		b"1111110100100101111110",
		b"1111110100010001110011",
		b"1111110011111110000110",
		b"1111110011101010111001",
		b"1111110011011000001100",
		b"1111110011000101111111",
		b"1111110010110100010100",
		b"1111110010100011001010",
		b"1111110010010010100010",
		b"1111110010000010011101",
		b"1111110001110010111011",
		b"1111110001100011111101",
		b"1111110001010101100011",
		b"1111110001000111101101",
		b"1111110000111010011101",
		b"1111110000101101110001",
		b"1111110000100001101011",
		b"1111110000010110001010",
		b"1111110000001011010000",
		b"1111110000000000111101",
		b"1111101111110111010000",
		b"1111101111101110001010",
		b"1111101111100101101011",
		b"1111101111011101110011",
		b"1111101111010110100011",
		b"1111101111001111111011",
		b"1111101111001001111010",
		b"1111101111000100100010",
		b"1111101110111111110001",
		b"1111101110111011101000",
		b"1111101110111000000111",
		b"1111101110110101001110",
		b"1111101110110010111101",
		b"1111101110110001010101",
		b"1111101110110000010100",
		b"1111101110101111111011",
		b"1111101110110000001001",
		b"1111101110110000111111",
		b"1111101110110010011101",
		b"1111101110110100100010",
		b"1111101110110111001110",
		b"1111101110111010100001",
		b"1111101110111110011011",
		b"1111101111000010111011",
		b"1111101111001000000001",
		b"1111101111001101101101",
		b"1111101111010011111111",
		b"1111101111011010110101",
		b"1111101111100010010001",
		b"1111101111101010010001",
		b"1111101111110010110101",
		b"1111101111111011111101",
		b"1111110000000101101000",
		b"1111110000001111110101",
		b"1111110000011010100101",
		b"1111110000100101110111",
		b"1111110000110001101010",
		b"1111110000111101111110",
		b"1111110001001010110010",
		b"1111110001011000000110",
		b"1111110001100101111001",
		b"1111110001110100001011",
		b"1111110010000010111010",
		b"1111110010010010000111",
		b"1111110010100001110000",
		b"1111110010110001110110",
		b"1111110011000010010111",
		b"1111110011010011010010",
		b"1111110011100100101000",
		b"1111110011110110010111",
		b"1111110100001000011111",
		b"1111110100011010111110",
		b"1111110100101101110101",
		b"1111110101000001000010",
		b"1111110101010100100101",
		b"1111110101101000011100",
		b"1111110101111100101000",
		b"1111110110010001001000",
		b"1111110110100101111001",
		b"1111110110111010111101",
		b"1111110111010000010001",
		b"1111110111100101110110",
		b"1111110111111011101010",
		b"1111111000010001101101",
		b"1111111000100111111101",
		b"1111111000111110011010",
		b"1111111001010101000011",
		b"1111111001101011110111",
		b"1111111010000010110101",
		b"1111111010011001111101",
		b"1111111010110001001101",
		b"1111111011001000100110",
		b"1111111011100000000101",
		b"1111111011110111101010",
		b"1111111100001111010100",
		b"1111111100100111000010",
		b"1111111100111110110100",
		b"1111111101010110101001",
		b"1111111101101110011111",
		b"1111111110000110010110",
		b"1111111110011110001101",
		b"1111111110110110000011",
		b"1111111111001101110111",
		b"1111111111100101101001",
		b"1111111111111101010111",
		b"0000000000010101000001",
		b"0000000000101100100110",
		b"0000000001000100000101",
		b"0000000001011011011101",
		b"0000000001110010101110",
		b"0000000010001001110110",
		b"0000000010100000110101",
		b"0000000010110111101010",
		b"0000000011001110010100",
		b"0000000011100100110011",
		b"0000000011111011000101",
		b"0000000100010001001011",
		b"0000000100100111000010",
		b"0000000100111100101011",
		b"0000000101010010000100",
		b"0000000101100111001110",
		b"0000000101111100000111",
		b"0000000110010000101110",
		b"0000000110100101000011",
		b"0000000110111001000101",
		b"0000000111001100110100",
		b"0000000111100000001110",
		b"0000000111110011010100",
		b"0000001000000110000101",
		b"0000001000011000011111",
		b"0000001000101010100011",
		b"0000001000111100001111",
		b"0000001001001101100100",
		b"0000001001011110100001",
		b"0000001001101111000100",
		b"0000001001111111001110",
		b"0000001010001110111111",
		b"0000001010011110010101",
		b"0000001010101101010000",
		b"0000001010111011110000",
		b"0000001011001001110100",
		b"0000001011010111011100",
		b"0000001011100100100111",
		b"0000001011110001010101",
		b"0000001011111101100110",
		b"0000001100001001011001",
		b"0000001100010100101111",
		b"0000001100011111100110",
		b"0000001100101001111110",
		b"0000001100110011110111",
		b"0000001100111101010001",
		b"0000001101000110001100",
		b"0000001101001110100110",
		b"0000001101010110100001",
		b"0000001101011101111100",
		b"0000001101100100110111",
		b"0000001101101011010001",
		b"0000001101110001001011",
		b"0000001101110110100011",
		b"0000001101111011011100",
		b"0000001101111111110011",
		b"0000001110000011101001",
		b"0000001110000110111110",
		b"0000001110001001110011",
		b"0000001110001100000110",
		b"0000001110001101111000",
		b"0000001110001111001010",
		b"0000001110001111111010",
		b"0000001110010000001010",
		b"0000001110001111111001",
		b"0000001110001111000111",
		b"0000001110001101110101",
		b"0000001110001100000010",
		b"0000001110001001101111",
		b"0000001110000110111100",
		b"0000001110000011101001",
		b"0000001101111111110110",
		b"0000001101111011100100",
		b"0000001101110110110011",
		b"0000001101110001100010",
		b"0000001101101011110011",
		b"0000001101100101100110",
		b"0000001101011110111011",
		b"0000001101010111110010",
		b"0000001101010000001011",
		b"0000001101001000000111",
		b"0000001100111111100111",
		b"0000001100110110101011",
		b"0000001100101101010010",
		b"0000001100100011011110",
		b"0000001100011001001111",
		b"0000001100001110100110",
		b"0000001100000011100010",
		b"0000001011111000000100",
		b"0000001011101100001110",
		b"0000001011011111111110",
		b"0000001011010011010111",
		b"0000001011000110011000",
		b"0000001010111001000001",
		b"0000001010101011010100",
		b"0000001010011101010010",
		b"0000001010001110111001",
		b"0000001010000000001100",
		b"0000001001110001001010",
		b"0000001001100001110101",
		b"0000001001010010001100",
		b"0000001001000010010001",
		b"0000001000110010000100",
		b"0000001000100001100110",
		b"0000001000010000111000",
		b"0000000111111111111001",
		b"0000000111101110101011",
		b"0000000111011101001110",
		b"0000000111001011100100",
		b"0000000110111001101100",
		b"0000000110100111100111",
		b"0000000110010101010111",
		b"0000000110000010111011",
		b"0000000101110000010101",
		b"0000000101011101100101",
		b"0000000101001010101011",
		b"0000000100110111101001",
		b"0000000100100100100000",
		b"0000000100010001001111",
		b"0000000011111101111000",
		b"0000000011101010011100",
		b"0000000011010110111010",
		b"0000000011000011010100",
		b"0000000010101111101011",
		b"0000000010011011111111",
		b"0000000010001000010001",
		b"0000000001110100100010",
		b"0000000001100000110001",
		b"0000000001001101000001",
		b"0000000000111001010010",
		b"0000000000100101100100",
		b"0000000000010001111001",
		b"1111111111111110010000",
		b"1111111111101010101011",
		b"1111111111010111001010",
		b"1111111111000011101110",
		b"1111111110110000011000",
		b"1111111110011101001000",
		b"1111111110001001111111",
		b"1111111101110110111110",
		b"1111111101100100000100",
		b"1111111101010001010100",
		b"1111111100111110101110",
		b"1111111100101100010010",
		b"1111111100011010000000",
		b"1111111100000111111011",
		b"1111111011110110000001",
		b"1111111011100100010100",
		b"1111111011010010110100",
		b"1111111011000001100010",
		b"1111111010110000011111",
		b"1111111010011111101011",
		b"1111111010001111000110",
		b"1111111001111110110010",
		b"1111111001101110101110",
		b"1111111001011110111100",
		b"1111111001001111011011",
		b"1111111001000000001101",
		b"1111111000110001010001",
		b"1111111000100010101001",
		b"1111111000010100010100",
		b"1111111000000110010100",
		b"1111110111111000101000",
		b"1111110111101011010001",
		b"1111110111011110010000",
		b"1111110111010001100100",
		b"1111110111000101001111",
		b"1111110110111001010000",
		b"1111110110101101101001",
		b"1111110110100010011001",
		b"1111110110010111100000",
		b"1111110110001101000000",
		b"1111110110000010111000",
		b"1111110101111001001000",
		b"1111110101101111110001",
		b"1111110101100110110100",
		b"1111110101011110010000",
		b"1111110101010110000110",
		b"1111110101001110010101",
		b"1111110101000110111111",
		b"1111110101000000000011",
		b"1111110100111001100001",
		b"1111110100110011011010",
		b"1111110100101101101110",
		b"1111110100101000011101",
		b"1111110100100011100110",
		b"1111110100011111001011",
		b"1111110100011011001011",
		b"1111110100010111100110",
		b"1111110100010100011101",
		b"1111110100010001101110",
		b"1111110100001111011100",
		b"1111110100001101100100",
		b"1111110100001100001000",
		b"1111110100001011000111",
		b"1111110100001010100010",
		b"1111110100001010010111",
		b"1111110100001010101000",
		b"1111110100001011010100",
		b"1111110100001100011011",
		b"1111110100001101111101",
		b"1111110100001111111010",
		b"1111110100010010010001",
		b"1111110100010101000011",
		b"1111110100011000001111",
		b"1111110100011011110101",
		b"1111110100011111110100",
		b"1111110100100100001110",
		b"1111110100101001000001",
		b"1111110100101110001101",
		b"1111110100110011110010",
		b"1111110100111001110000",
		b"1111110101000000000110",
		b"1111110101000110110100",
		b"1111110101001101111010",
		b"1111110101010101010111",
		b"1111110101011101001100",
		b"1111110101100101010111",
		b"1111110101101101111001",
		b"1111110101110110110001",
		b"1111110101111111111110",
		b"1111110110001001100001",
		b"1111110110010011011001",
		b"1111110110011101100101",
		b"1111110110101000000101",
		b"1111110110110010111001",
		b"1111110110111110000000",
		b"1111110111001001011010",
		b"1111110111010101000101",
		b"1111110111100001000011",
		b"1111110111101101010010",
		b"1111110111111001110010",
		b"1111111000000110100011",
		b"1111111000010011100011",
		b"1111111000100000110010",
		b"1111111000101110010001",
		b"1111111000111011111101",
		b"1111111001001001110111",
		b"1111111001010111111111",
		b"1111111001100110010011",
		b"1111111001110100110100",
		b"1111111010000011100000",
		b"1111111010010010010111",
		b"1111111010100001011000",
		b"1111111010110000100100",
		b"1111111010111111111000",
		b"1111111011001111010110",
		b"1111111011011110111011",
		b"1111111011101110101000",
		b"1111111011111110011101",
		b"1111111100001110010111",
		b"1111111100011110011000",
		b"1111111100101110011101",
		b"1111111100111110101000",
		b"1111111101001110110110",
		b"1111111101011111001000",
		b"1111111101101111011101",
		b"1111111101111111110100",
		b"1111111110010000001101",
		b"1111111110100000100111",
		b"1111111110110001000001",
		b"1111111111000001011100",
		b"1111111111010001110101",
		b"1111111111100010001110",
		b"1111111111110010100100",
		b"0000000000000010111000",
		b"0000000000010011001010",
		b"0000000000100011010111",
		b"0000000000110011100001",
		b"0000000001000011100110",
		b"0000000001010011100101",
		b"0000000001100011011111",
		b"0000000001110011010010",
		b"0000000010000010111111",
		b"0000000010010010100100",
		b"0000000010100010000001",
		b"0000000010110001010101",
		b"0000000011000000100001",
		b"0000000011001111100011",
		b"0000000011011110011011",
		b"0000000011101101001000",
		b"0000000011111011101010",
		b"0000000100001010000000",
		b"0000000100011000001011",
		b"0000000100100110001001",
		b"0000000100110011111010",
		b"0000000101000001011101",
		b"0000000101001110110011",
		b"0000000101011011111010",
		b"0000000101101000110011",
		b"0000000101110101011100",
		b"0000000110000001110110",
		b"0000000110001110000000",
		b"0000000110011001111001",
		b"0000000110100101100010",
		b"0000000110110000111010",
		b"0000000110111100000000",
		b"0000000111000110110100",
		b"0000000111010001010110",
		b"0000000111011011100101",
		b"0000000111100101100010",
		b"0000000111101111001011",
		b"0000000111111000100010",
		b"0000001000000001100100",
		b"0000001000001010010010",
		b"0000001000010010101101",
		b"0000001000011010110011",
		b"0000001000100010100100",
		b"0000001000101010000000",
		b"0000001000110001000111",
		b"0000001000110111111000",
		b"0000001000111110010101",
		b"0000001001000100011011",
		b"0000001001001010001100",
		b"0000001001001111100111",
		b"0000001001010100101011",
		b"0000001001011001011001",
		b"0000001001011101110001",
		b"0000001001100001110011",
		b"0000001001100101011110",
		b"0000001001101000110011",
		b"0000001001101011110000",
		b"0000001001101110010111",
		b"0000001001110000101000",
		b"0000001001110010100010",
		b"0000001001110100000100",
		b"0000001001110101010001",
		b"0000001001110110000110",
		b"0000001001110110100101",
		b"0000001001110110101101",
		b"0000001001110110011111",
		b"0000001001110101111010",
		b"0000001001110100111110",
		b"0000001001110011101101",
		b"0000001001110010000101",
		b"0000001001110000000111",
		b"0000001001101101110011",
		b"0000001001101011001001",
		b"0000001001101000001010",
		b"0000001001100100110101",
		b"0000001001100001001010",
		b"0000001001011101001011",
		b"0000001001011000110111",
		b"0000001001010100001101",
		b"0000001001001111010000",
		b"0000001001001001111110",
		b"0000001001000100011000",
		b"0000001000111110011111",
		b"0000001000111000010001",
		b"0000001000110001110001",
		b"0000001000101010111110",
		b"0000001000100011111000",
		b"0000001000011100100000",
		b"0000001000010100110101",
		b"0000001000001100111001",
		b"0000001000000100101100",
		b"0000000111111100001110",
		b"0000000111110011011110",
		b"0000000111101010011111",
		b"0000000111100001010000",
		b"0000000111010111110001",
		b"0000000111001110000011",
		b"0000000111000100000110",
		b"0000000110111001111011",
		b"0000000110101111100001",
		b"0000000110100100111010",
		b"0000000110011010000110",
		b"0000000110001111000110",
		b"0000000110000011111000",
		b"0000000101111000011111",
		b"0000000101101100111011",
		b"0000000101100001001011",
		b"0000000101010101010001",
		b"0000000101001001001101",
		b"0000000100111101000000",
		b"0000000100110000101001",
		b"0000000100100100001001",
		b"0000000100010111100001",
		b"0000000100001010110001",
		b"0000000011111101111011",
		b"0000000011110000111101",
		b"0000000011100011111001",
		b"0000000011010110101111",
		b"0000000011001001100000",
		b"0000000010111100001011",
		b"0000000010101110110011",
		b"0000000010100001010110",
		b"0000000010010011110111",
		b"0000000010000110010100",
		b"0000000001111000101111",
		b"0000000001101011001000",
		b"0000000001011101011111",
		b"0000000001001111110110",
		b"0000000001000010001100",
		b"0000000000110100100010",
		b"0000000000100110111001",
		b"0000000000011001010001",
		b"0000000000001011101010",
		b"1111111111111110000101",
		b"1111111111110000100011",
		b"1111111111100011000100",
		b"1111111111010101101000",
		b"1111111111001000010000",
		b"1111111110111010111100",
		b"1111111110101101101101",
		b"1111111110100000100011",
		b"1111111110010011011111",
		b"1111111110000110100010",
		b"1111111101111001101011",
		b"1111111101101100111011",
		b"1111111101100000010010",
		b"1111111101010011110001",
		b"1111111101000111011001",
		b"1111111100111011001010",
		b"1111111100101111000011",
		b"1111111100100011000111",
		b"1111111100010111010100",
		b"1111111100001011101100",
		b"1111111100000000001110",
		b"1111111011110100111100",
		b"1111111011101001110101",
		b"1111111011011110111010",
		b"1111111011010100001011",
		b"1111111011001001101001",
		b"1111111010111111010100",
		b"1111111010110101001100",
		b"1111111010101011010010",
		b"1111111010100001100110",
		b"1111111010011000000111",
		b"1111111010001110111000",
		b"1111111010000101110111",
		b"1111111001111101000101",
		b"1111111001110100100011",
		b"1111111001101100010000",
		b"1111111001100100001101",
		b"1111111001011100011011",
		b"1111111001010100111000",
		b"1111111001001101100110",
		b"1111111001000110100101",
		b"1111111000111111110101",
		b"1111111000111001010111",
		b"1111111000110011001001",
		b"1111111000101101001101",
		b"1111111000100111100011",
		b"1111111000100010001011",
		b"1111111000011101000100",
		b"1111111000011000010000",
		b"1111111000010011101110",
		b"1111111000001111011111",
		b"1111111000001011100010",
		b"1111111000000111110111",
		b"1111111000000100011111",
		b"1111111000000001011010",
		b"1111110111111110101000",
		b"1111110111111100001000",
		b"1111110111111001111011",
		b"1111110111111000000010",
		b"1111110111110110011011",
		b"1111110111110101000110",
		b"1111110111110100000101",
		b"1111110111110011010111",
		b"1111110111110010111100",
		b"1111110111110010110011",
		b"1111110111110010111101",
		b"1111110111110011011010",
		b"1111110111110100001001",
		b"1111110111110101001011",
		b"1111110111110110100000",
		b"1111110111111000000111",
		b"1111110111111010000000",
		b"1111110111111100001011",
		b"1111110111111110101000",
		b"1111111000000001011000",
		b"1111111000000100011001",
		b"1111111000000111101011",
		b"1111111000001011001111",
		b"1111111000001111000100",
		b"1111111000010011001010",
		b"1111111000010111100001",
		b"1111111000011100001001",
		b"1111111000100001000001",
		b"1111111000100110001001",
		b"1111111000101011100010",
		b"1111111000110001001010",
		b"1111111000110111000010",
		b"1111111000111101001000",
		b"1111111001000011011110",
		b"1111111001001010000011",
		b"1111111001010000110110",
		b"1111111001010111110111",
		b"1111111001011111000110",
		b"1111111001100110100011",
		b"1111111001101110001101",
		b"1111111001110110000100",
		b"1111111001111110000111",
		b"1111111010000110010111",
		b"1111111010001110110011",
		b"1111111010010111011011",
		b"1111111010100000001110",
		b"1111111010101001001100",
		b"1111111010110010010100",
		b"1111111010111011100111",
		b"1111111011000101000100",
		b"1111111011001110101010",
		b"1111111011011000011010",
		b"1111111011100010010010",
		b"1111111011101100010011",
		b"1111111011110110011100",
		b"1111111100000000101100",
		b"1111111100001011000100",
		b"1111111100010101100010",
		b"1111111100100000000111",
		b"1111111100101010110011",
		b"1111111100110101100100",
		b"1111111101000000011010",
		b"1111111101001011010101",
		b"1111111101010110010100",
		b"1111111101100001011000",
		b"1111111101101100100000",
		b"1111111101110111101010",
		b"1111111110000010111000",
		b"1111111110001110001000",
		b"1111111110011001011010",
		b"1111111110100100101110",
		b"1111111110110000000011",
		b"1111111110111011011000",
		b"1111111111000110101111",
		b"1111111111010010000101",
		b"1111111111011101011011",
		b"1111111111101000110000",
		b"1111111111110100000100",
		b"1111111111111111010110",
		b"0000000000001010100110",
		b"0000000000010101110100",
		b"0000000000100000111111",
		b"0000000000101100000111",
		b"0000000000110111001100",
		b"0000000001000010001100",
		b"0000000001001101001000",
		b"0000000001011000000000",
		b"0000000001100010110010",
		b"0000000001101101011111",
		b"0000000001111000000110",
		b"0000000010000010100111",
		b"0000000010001101000010",
		b"0000000010010111010101",
		b"0000000010100001100001",
		b"0000000010101011100110",
		b"0000000010110101100011",
		b"0000000010111111011000",
		b"0000000011001001000100",
		b"0000000011010010100111",
		b"0000000011011100000001",
		b"0000000011100101010001",
		b"0000000011101110011000",
		b"0000000011110111010100",
		b"0000000100000000000110",
		b"0000000100001000101101",
		b"0000000100010001001010",
		b"0000000100011001011011",
		b"0000000100100001100000",
		b"0000000100101001011010",
		b"0000000100110001001000",
		b"0000000100111000101010",
		b"0000000100111111111111",
		b"0000000101000111000111",
		b"0000000101001110000011",
		b"0000000101010100110001",
		b"0000000101011011010010",
		b"0000000101100001100101",
		b"0000000101100111101011",
		b"0000000101101101100011",
		b"0000000101110011001101",
		b"0000000101111000101000",
		b"0000000101111101110101",
		b"0000000110000010110100",
		b"0000000110000111100100",
		b"0000000110001100000101",
		b"0000000110010000010111",
		b"0000000110010100011011",
		b"0000000110011000001111",
		b"0000000110011011110011",
		b"0000000110011111001001",
		b"0000000110100010001111",
		b"0000000110100101000110",
		b"0000000110100111101101",
		b"0000000110101010000101",
		b"0000000110101100001101",
		b"0000000110101110000101",
		b"0000000110101111101110",
		b"0000000110110001000111",
		b"0000000110110010010000",
		b"0000000110110011001010",
		b"0000000110110011110100",
		b"0000000110110100001110",
		b"0000000110110100011001",
		b"0000000110110100010101",
		b"0000000110110100000000",
		b"0000000110110011011101",
		b"0000000110110010101001",
		b"0000000110110001100111",
		b"0000000110110000010101",
		b"0000000110101110110100",
		b"0000000110101101000100",
		b"0000000110101011000101",
		b"0000000110101000111000",
		b"0000000110100110011011",
		b"0000000110100011110000",
		b"0000000110100000110110",
		b"0000000110011101101111",
		b"0000000110011010011001",
		b"0000000110010110110100",
		b"0000000110010011000011",
		b"0000000110001111000011",
		b"0000000110001010110110",
		b"0000000110000110011100",
		b"0000000110000001110100",
		b"0000000101111101000000",
		b"0000000101110111111111",
		b"0000000101110010110001",
		b"0000000101101101010111",
		b"0000000101100111110001",
		b"0000000101100010000000",
		b"0000000101011100000010",
		b"0000000101010101111010",
		b"0000000101001111100110",
		b"0000000101001001001000",
		b"0000000101000010011111",
		b"0000000100111011101100",
		b"0000000100110100101110",
		b"0000000100101101100111",
		b"0000000100100110010111",
		b"0000000100011110111101",
		b"0000000100010111011011",
		b"0000000100001111110000",
		b"0000000100000111111100",
		b"0000000100000000000001",
		b"0000000011110111111110",
		b"0000000011101111110100",
		b"0000000011100111100010",
		b"0000000011011111001010",
		b"0000000011010110101011",
		b"0000000011001110000110",
		b"0000000011000101011100",
		b"0000000010111100101100",
		b"0000000010110011110111",
		b"0000000010101010111101",
		b"0000000010100001111110",
		b"0000000010011000111100",
		b"0000000010001111110101",
		b"0000000010000110101011",
		b"0000000001111101011110",
		b"0000000001110100001111",
		b"0000000001101010111100",
		b"0000000001100001101000",
		b"0000000001011000010010",
		b"0000000001001110111010",
		b"0000000001000101100001",
		b"0000000000111100000111",
		b"0000000000110010101101",
		b"0000000000101001010011",
		b"0000000000011111111001",
		b"0000000000010110100000",
		b"0000000000001101001000",
		b"0000000000000011110000",
		b"1111111111111010011011",
		b"1111111111110001000111",
		b"1111111111100111110101",
		b"1111111111011110100110",
		b"1111111111010101011010",
		b"1111111111001100010001",
		b"1111111111000011001100",
		b"1111111110111010001010",
		b"1111111110110001001100",
		b"1111111110101000010011",
		b"1111111110011111011111",
		b"1111111110010110101111",
		b"1111111110001110000101",
		b"1111111110000101100001",
		b"1111111101111101000010",
		b"1111111101110100101010",
		b"1111111101101100011000",
		b"1111111101100100001100",
		b"1111111101011100001000",
		b"1111111101010100001011",
		b"1111111101001100010110",
		b"1111111101000100101000",
		b"1111111100111101000011",
		b"1111111100110101100110",
		b"1111111100101110010001",
		b"1111111100100111000101",
		b"1111111100100000000010",
		b"1111111100011001001001",
		b"1111111100010010011000",
		b"1111111100001011110010",
		b"1111111100000101010101",
		b"1111111011111111000011",
		b"1111111011111000111010",
		b"1111111011110010111100",
		b"1111111011101101001001",
		b"1111111011100111100001",
		b"1111111011100010000011",
		b"1111111011011100110001",
		b"1111111011010111101010",
		b"1111111011010010101111",
		b"1111111011001101111111",
		b"1111111011001001011010",
		b"1111111011000101000010",
		b"1111111011000000110110",
		b"1111111010111100110110",
		b"1111111010111001000001",
		b"1111111010110101011010",
		b"1111111010110001111110",
		b"1111111010101110110000",
		b"1111111010101011101101",
		b"1111111010101000111000",
		b"1111111010100110001111",
		b"1111111010100011110010",
		b"1111111010100001100011",
		b"1111111010011111100000",
		b"1111111010011101101011",
		b"1111111010011100000010",
		b"1111111010011010100110",
		b"1111111010011001010111",
		b"1111111010011000010101",
		b"1111111010010111100000",
		b"1111111010010110111000",
		b"1111111010010110011101",
		b"1111111010010110001111",
		b"1111111010010110001110",
		b"1111111010010110011001",
		b"1111111010010110110010",
		b"1111111010010111010111",
		b"1111111010011000001001",
		b"1111111010011001000111",
		b"1111111010011010010010",
		b"1111111010011011101010",
		b"1111111010011101001101",
		b"1111111010011110111110",
		b"1111111010100000111010",
		b"1111111010100011000010",
		b"1111111010100101010111",
		b"1111111010100111110111",
		b"1111111010101010100011",
		b"1111111010101101011011",
		b"1111111010110000011110",
		b"1111111010110011101101",
		b"1111111010110111000111",
		b"1111111010111010101011",
		b"1111111010111110011011",
		b"1111111011000010010101",
		b"1111111011000110011010",
		b"1111111011001010101010",
		b"1111111011001111000011",
		b"1111111011010011100111",
		b"1111111011011000010100",
		b"1111111011011101001011",
		b"1111111011100010001100",
		b"1111111011100111010101",
		b"1111111011101100101000",
		b"1111111011110010000011",
		b"1111111011110111100111",
		b"1111111011111101010100",
		b"1111111100000011001000",
		b"1111111100001001000101",
		b"1111111100001111001001",
		b"1111111100010101010100",
		b"1111111100011011100111",
		b"1111111100100010000000",
		b"1111111100101000100001",
		b"1111111100101111000111",
		b"1111111100110101110100",
		b"1111111100111100100111",
		b"1111111101000011100000",
		b"1111111101001010011110",
		b"1111111101010001100001",
		b"1111111101011000101001",
		b"1111111101011111110101",
		b"1111111101100111000110",
		b"1111111101101110011011",
		b"1111111101110101110100",
		b"1111111101111101010001",
		b"1111111110000100110000",
		b"1111111110001100010011",
		b"1111111110010011111000",
		b"1111111110011011100000",
		b"1111111110100011001010",
		b"1111111110101010110110",
		b"1111111110110010100011",
		b"1111111110111010010010",
		b"1111111111000010000010",
		b"1111111111001001110010",
		b"1111111111010001100011",
		b"1111111111011001010101",
		b"1111111111100001000110",
		b"1111111111101000110111",
		b"1111111111110000100111",
		b"1111111111111000010110",
		b"0000000000000000000100",
		b"0000000000000111110001",
		b"0000000000001111011100",
		b"0000000000010111000101",
		b"0000000000011110101100",
		b"0000000000100110010000",
		b"0000000000101101110001",
		b"0000000000110101010000",
		b"0000000000111100101011",
		b"0000000001000100000011",
		b"0000000001001011010111",
		b"0000000001010010100111",
		b"0000000001011001110010",
		b"0000000001100000111001",
		b"0000000001100111111100",
		b"0000000001101110111001",
		b"0000000001110101110001",
		b"0000000001111100100100",
		b"0000000010000011010001",
		b"0000000010001001111000",
		b"0000000010010000011001",
		b"0000000010010110110100",
		b"0000000010011101001000",
		b"0000000010100011010101",
		b"0000000010101001011100",
		b"0000000010101111011011",
		b"0000000010110101010011",
		b"0000000010111011000011",
		b"0000000011000000101100",
		b"0000000011000110001101",
		b"0000000011001011100110",
		b"0000000011010000110110",
		b"0000000011010101111110",
		b"0000000011011010111110",
		b"0000000011011111110101",
		b"0000000011100100100011",
		b"0000000011101001001000",
		b"0000000011101101100100",
		b"0000000011110001110111",
		b"0000000011110110000000",
		b"0000000011111010000000",
		b"0000000011111101110111",
		b"0000000100000001100011",
		b"0000000100000101000110",
		b"0000000100001000011111",
		b"0000000100001011101110",
		b"0000000100001110110011",
		b"0000000100010001101101",
		b"0000000100010100011101",
		b"0000000100010111000100",
		b"0000000100011001011111",
		b"0000000100011011110000",
		b"0000000100011101110111",
		b"0000000100011111110100",
		b"0000000100100001100101",
		b"0000000100100011001100",
		b"0000000100100100101001",
		b"0000000100100101111011",
		b"0000000100100111000010",
		b"0000000100100111111110",
		b"0000000100101000110000",
		b"0000000100101001011000",
		b"0000000100101001110100",
		b"0000000100101010000110",
		b"0000000100101010001101",
		b"0000000100101010001010",
		b"0000000100101001111100",
		b"0000000100101001100100",
		b"0000000100101001000001",
		b"0000000100101000010100",
		b"0000000100100111011100",
		b"0000000100100110011011",
		b"0000000100100101001111",
		b"0000000100100011111000",
		b"0000000100100010011000",
		b"0000000100100000101110",
		b"0000000100011110111001",
		b"0000000100011100111011",
		b"0000000100011010110011",
		b"0000000100011000100010",
		b"0000000100010110000111",
		b"0000000100010011100011",
		b"0000000100010000110101",
		b"0000000100001101111110",
		b"0000000100001010111111",
		b"0000000100000111110110",
		b"0000000100000100100101",
		b"0000000100000001001011",
		b"0000000011111101101000",
		b"0000000011111001111101",
		b"0000000011110110001010",
		b"0000000011110010001111",
		b"0000000011101110001101",
		b"0000000011101010000010",
		b"0000000011100101110000",
		b"0000000011100001010111",
		b"0000000011011100110110",
		b"0000000011011000001111",
		b"0000000011010011100001",
		b"0000000011001110101100",
		b"0000000011001001110001",
		b"0000000011000100101111",
		b"0000000010111111101000",
		b"0000000010111010011010",
		b"0000000010110101000111",
		b"0000000010101111101111",
		b"0000000010101010010010",
		b"0000000010100100101111",
		b"0000000010011111001000",
		b"0000000010011001011100",
		b"0000000010010011101100",
		b"0000000010001101110111",
		b"0000000010000111111111",
		b"0000000010000010000011",
		b"0000000001111100000011",
		b"0000000001110110000000",
		b"0000000001101111111011",
		b"0000000001101001110010",
		b"0000000001100011100111",
		b"0000000001011101011001",
		b"0000000001010111001001",
		b"0000000001010000111000",
		b"0000000001001010100100",
		b"0000000001000100010000",
		b"0000000000111101111010",
		b"0000000000110111100011",
		b"0000000000110001001011",
		b"0000000000101010110011",
		b"0000000000100100011010",
		b"0000000000011110000001",
		b"0000000000010111101001",
		b"0000000000010001010001",
		b"0000000000001010111001",
		b"0000000000000100100010",
		b"1111111111111110001100",
		b"1111111111110111111000",
		b"1111111111110001100101",
		b"1111111111101011010011",
		b"1111111111100101000100",
		b"1111111111011110110111",
		b"1111111111011000101100",
		b"1111111111010010100011",
		b"1111111111001100011110",
		b"1111111111000110011011",
		b"1111111111000000011011",
		b"1111111110111010011111",
		b"1111111110110100100111",
		b"1111111110101110110010",
		b"1111111110101001000001",
		b"1111111110100011010100",
		b"1111111110011101101100",
		b"1111111110011000001000",
		b"1111111110010010101001",
		b"1111111110001101001111",
		b"1111111110000111111010",
		b"1111111110000010101010",
		b"1111111101111101011111",
		b"1111111101111000011011",
		b"1111111101110011011011",
		b"1111111101101110100010",
		b"1111111101101001101111",
		b"1111111101100101000010",
		b"1111111101100000011011",
		b"1111111101011011111011",
		b"1111111101010111100010",
		b"1111111101010011001111",
		b"1111111101001111000011",
		b"1111111101001010111111",
		b"1111111101000111000001",
		b"1111111101000011001011",
		b"1111111100111111011100",
		b"1111111100111011110100",
		b"1111111100111000010100",
		b"1111111100110100111100",
		b"1111111100110001101100",
		b"1111111100101110100100",
		b"1111111100101011100011",
		b"1111111100101000101011",
		b"1111111100100101111011",
		b"1111111100100011010010",
		b"1111111100100000110011",
		b"1111111100011110011011",
		b"1111111100011100001100",
		b"1111111100011010000110",
		b"1111111100011000001000",
		b"1111111100010110010010",
		b"1111111100010100100101",
		b"1111111100010011000001",
		b"1111111100010001100101",
		b"1111111100010000010010",
		b"1111111100001111001000",
		b"1111111100001110000110",
		b"1111111100001101001110",
		b"1111111100001100011101",
		b"1111111100001011110110",
		b"1111111100001011010111",
		b"1111111100001011000001",
		b"1111111100001010110100",
		b"1111111100001010101111",
		b"1111111100001010110011",
		b"1111111100001011000000",
		b"1111111100001011010101",
		b"1111111100001011110011",
		b"1111111100001100011001",
		b"1111111100001101001000",
		b"1111111100001101111111",
		b"1111111100001110111111",
		b"1111111100010000000111",
		b"1111111100010001010111",
		b"1111111100010010101111",
		b"1111111100010100001111",
		b"1111111100010101111000",
		b"1111111100010111101000",
		b"1111111100011001100000",
		b"1111111100011011100000",
		b"1111111100011101100111",
		b"1111111100011111110111",
		b"1111111100100010001101",
		b"1111111100100100101011",
		b"1111111100100111010000",
		b"1111111100101001111100",
		b"1111111100101100110000",
		b"1111111100101111101010",
		b"1111111100110010101011",
		b"1111111100110101110010",
		b"1111111100111001000000",
		b"1111111100111100010101",
		b"1111111100111111101111",
		b"1111111101000011010000",
		b"1111111101000110110111",
		b"1111111101001010100100",
		b"1111111101001110010110",
		b"1111111101010010001110",
		b"1111111101010110001011",
		b"1111111101011010001101",
		b"1111111101011110010100",
		b"1111111101100010100001",
		b"1111111101100110110010",
		b"1111111101101011000111",
		b"1111111101101111100001",
		b"1111111101110011111111",
		b"1111111101111000100010",
		b"1111111101111101001000",
		b"1111111110000001110001",
		b"1111111110000110011111",
		b"1111111110001011001111",
		b"1111111110010000000011",
		b"1111111110010100111010",
		b"1111111110011001110100",
		b"1111111110011110110000",
		b"1111111110100011101111",
		b"1111111110101000110000",
		b"1111111110101101110011",
		b"1111111110110010111000",
		b"1111111110110111111111",
		b"1111111110111101000111",
		b"1111111111000010010001",
		b"1111111111000111011011",
		b"1111111111001100100111",
		b"1111111111010001110100",
		b"1111111111010111000001",
		b"1111111111011100001110",
		b"1111111111100001011100",
		b"1111111111100110101010",
		b"1111111111101011111000",
		b"1111111111110001000101",
		b"1111111111110110010010",
		b"1111111111111011011110",
		b"0000000000000000101001",
		b"0000000000000101110011",
		b"0000000000001010111100",
		b"0000000000010000000100",
		b"0000000000010101001010",
		b"0000000000011010001110",
		b"0000000000011111010001",
		b"0000000000100100010001",
		b"0000000000101001001111",
		b"0000000000101110001011",
		b"0000000000110011000100",
		b"0000000000110111111010",
		b"0000000000111100101101",
		b"0000000001000001011101",
		b"0000000001000110001010",
		b"0000000001001010110100",
		b"0000000001001111011010",
		b"0000000001010011111100",
		b"0000000001011000011011",
		b"0000000001011100110101",
		b"0000000001100001001011",
		b"0000000001100101011101",
		b"0000000001101001101011",
		b"0000000001101101110100",
		b"0000000001110001111000",
		b"0000000001110101111000",
		b"0000000001111001110010",
		b"0000000001111101101000",
		b"0000000010000001011000",
		b"0000000010000101000011",
		b"0000000010001000101001",
		b"0000000010001100001001",
		b"0000000010001111100011",
		b"0000000010010010111000",
		b"0000000010010110000111",
		b"0000000010011001010000",
		b"0000000010011100010011",
		b"0000000010011111010000",
		b"0000000010100010000110",
		b"0000000010100100110111",
		b"0000000010100111100001",
		b"0000000010101010000100",
		b"0000000010101100100001",
		b"0000000010101110111000",
		b"0000000010110001001000",
		b"0000000010110011010001",
		b"0000000010110101010100",
		b"0000000010110111001111",
		b"0000000010111001000100",
		b"0000000010111010110010",
		b"0000000010111100011001",
		b"0000000010111101111001",
		b"0000000010111111010010",
		b"0000000011000000100101",
		b"0000000011000001110000",
		b"0000000011000010110100",
		b"0000000011000011110001",
		b"0000000011000100100110",
		b"0000000011000101010101",
		b"0000000011000101111101",
		b"0000000011000110011110",
		b"0000000011000110110111",
		b"0000000011000111001001",
		b"0000000011000111010101",
		b"0000000011000111011001",
		b"0000000011000111010110",
		b"0000000011000111001101",
		b"0000000011000110111100",
		b"0000000011000110100100",
		b"0000000011000110000110",
		b"0000000011000101100000",
		b"0000000011000100110100",
		b"0000000011000100000001",
		b"0000000011000011000111",
		b"0000000011000010000111",
		b"0000000011000000111111",
		b"0000000010111111110010",
		b"0000000010111110011110",
		b"0000000010111101000011",
		b"0000000010111011100010",
		b"0000000010111001111010",
		b"0000000010111000001101",
		b"0000000010110110011001",
		b"0000000010110100011111",
		b"0000000010110010100000",
		b"0000000010110000011010",
		b"0000000010101110001111",
		b"0000000010101011111101",
		b"0000000010101001100111",
		b"0000000010100111001011",
		b"0000000010100100101001",
		b"0000000010100010000010",
		b"0000000010011111010110",
		b"0000000010011100100101",
		b"0000000010011001101111",
		b"0000000010010110110100",
		b"0000000010010011110100",
		b"0000000010010000101111",
		b"0000000010001101100111",
		b"0000000010001010011001",
		b"0000000010000111001000",
		b"0000000010000011110011",
		b"0000000010000000011001",
		b"0000000001111100111100",
		b"0000000001111001011011",
		b"0000000001110101110110",
		b"0000000001110010001110",
		b"0000000001101110100011",
		b"0000000001101010110100",
		b"0000000001100111000011",
		b"0000000001100011001110",
		b"0000000001011111010111",
		b"0000000001011011011101",
		b"0000000001010111100001",
		b"0000000001010011100010",
		b"0000000001001111100010",
		b"0000000001001011011111",
		b"0000000001000111011011",
		b"0000000001000011010100",
		b"0000000000111111001101",
		b"0000000000111011000011",
		b"0000000000110110111001",
		b"0000000000110010101101",
		b"0000000000101110100001",
		b"0000000000101010010011",
		b"0000000000100110000101",
		b"0000000000100001110111",
		b"0000000000011101101000",
		b"0000000000011001011001",
		b"0000000000010101001010",
		b"0000000000010000111011",
		b"0000000000001100101100",
		b"0000000000001000011101",
		b"0000000000000100010000",
		b"0000000000000000000010",
		b"1111111111111011110110",
		b"1111111111110111101010",
		b"1111111111110011100000",
		b"1111111111101111010111",
		b"1111111111101011001111",
		b"1111111111100111001001",
		b"1111111111100011000101",
		b"1111111111011111000010",
		b"1111111111011011000001",
		b"1111111111010111000011",
		b"1111111111010011000110",
		b"1111111111001111001100",
		b"1111111111001011010100",
		b"1111111111000111011111",
		b"1111111111000011101101",
		b"1111111110111111111110",
		b"1111111110111100010001",
		b"1111111110111000101000",
		b"1111111110110101000010",
		b"1111111110110001011111",
		b"1111111110101101111111",
		b"1111111110101010100011",
		b"1111111110100111001011",
		b"1111111110100011110111",
		b"1111111110100000100110",
		b"1111111110011101011010",
		b"1111111110011010010001",
		b"1111111110010111001101",
		b"1111111110010100001101",
		b"1111111110010001010001",
		b"1111111110001110011010",
		b"1111111110001011100111",
		b"1111111110001000111001",
		b"1111111110000110001111",
		b"1111111110000011101011",
		b"1111111110000001001011",
		b"1111111101111110110000",
		b"1111111101111100011010",
		b"1111111101111010001001",
		b"1111111101110111111110",
		b"1111111101110101110111",
		b"1111111101110011110110",
		b"1111111101110001111010",
		b"1111111101110000000011",
		b"1111111101101110010010",
		b"1111111101101100100110",
		b"1111111101101010111111",
		b"1111111101101001011110",
		b"1111111101101000000011",
		b"1111111101100110101101",
		b"1111111101100101011101",
		b"1111111101100100010010",
		b"1111111101100011001101",
		b"1111111101100010001110",
		b"1111111101100001010101",
		b"1111111101100000100001",
		b"1111111101011111110011",
		b"1111111101011111001010",
		b"1111111101011110101000",
		b"1111111101011110001011",
		b"1111111101011101110011",
		b"1111111101011101100010",
		b"1111111101011101010110",
		b"1111111101011101010000",
		b"1111111101011101010000",
		b"1111111101011101010101",
		b"1111111101011101100000",
		b"1111111101011101110000",
		b"1111111101011110000110",
		b"1111111101011110100010",
		b"1111111101011111000011",
		b"1111111101011111101010",
		b"1111111101100000010110",
		b"1111111101100001000111",
		b"1111111101100001111110",
		b"1111111101100010111010",
		b"1111111101100011111100",
		b"1111111101100101000010",
		b"1111111101100110001110",
		b"1111111101100111011111",
		b"1111111101101000110101",
		b"1111111101101010010000",
		b"1111111101101011110000",
		b"1111111101101101010100",
		b"1111111101101110111110",
		b"1111111101110000101100",
		b"1111111101110010011111",
		b"1111111101110100010110",
		b"1111111101110110010010",
		b"1111111101111000010010",
		b"1111111101111010010111",
		b"1111111101111100011111",
		b"1111111101111110101100",
		b"1111111110000000111101",
		b"1111111110000011010010",
		b"1111111110000101101010",
		b"1111111110001000000111",
		b"1111111110001010100111",
		b"1111111110001101001010",
		b"1111111110001111110001",
		b"1111111110010010011100",
		b"1111111110010101001001",
		b"1111111110010111111010",
		b"1111111110011010101110",
		b"1111111110011101100100",
		b"1111111110100000011110",
		b"1111111110100011011010",
		b"1111111110100110011001",
		b"1111111110101001011010",
		b"1111111110101100011110",
		b"1111111110101111100100",
		b"1111111110110010101100",
		b"1111111110110101110110",
		b"1111111110111001000010",
		b"1111111110111100010000",
		b"1111111110111111011111",
		b"1111111111000010110000",
		b"1111111111000110000011",
		b"1111111111001001010110",
		b"1111111111001100101011",
		b"1111111111010000000001",
		b"1111111111010011011000",
		b"1111111111010110110000",
		b"1111111111011010001000",
		b"1111111111011101100001",
		b"1111111111100000111011",
		b"1111111111100100010101",
		b"1111111111100111101111",
		b"1111111111101011001001",
		b"1111111111101110100011",
		b"1111111111110001111101",
		b"1111111111110101010111",
		b"1111111111111000110001",
		b"1111111111111100001010",
		b"1111111111111111100010",
		b"0000000000000010111001",
		b"0000000000000110010000",
		b"0000000000001001100110",
		b"0000000000001100111011",
		b"0000000000010000001111",
		b"0000000000010011100001",
		b"0000000000010110110010",
		b"0000000000011010000001",
		b"0000000000011101001111",
		b"0000000000100000011011",
		b"0000000000100011100101",
		b"0000000000100110101110",
		b"0000000000101001110100",
		b"0000000000101100111000",
		b"0000000000101111111010",
		b"0000000000110010111010",
		b"0000000000110101110111",
		b"0000000000111000110001",
		b"0000000000111011101001",
		b"0000000000111110011111",
		b"0000000001000001010001",
		b"0000000001000100000001",
		b"0000000001000110101101",
		b"0000000001001001010111",
		b"0000000001001011111101",
		b"0000000001001110100001",
		b"0000000001010001000001",
		b"0000000001010011011101",
		b"0000000001010101110110",
		b"0000000001011000001100",
		b"0000000001011010011110",
		b"0000000001011100101100",
		b"0000000001011110110110",
		b"0000000001100000111101",
		b"0000000001100011000000",
		b"0000000001100100111111",
		b"0000000001100110111010",
		b"0000000001101000110001",
		b"0000000001101010100100",
		b"0000000001101100010011",
		b"0000000001101101111110",
		b"0000000001101111100100",
		b"0000000001110001000110",
		b"0000000001110010100100",
		b"0000000001110011111110",
		b"0000000001110101010011",
		b"0000000001110110100100",
		b"0000000001110111110000",
		b"0000000001111000111000",
		b"0000000001111001111011",
		b"0000000001111010111010",
		b"0000000001111011110101",
		b"0000000001111100101010",
		b"0000000001111101011100",
		b"0000000001111110001001",
		b"0000000001111110110001",
		b"0000000001111111010100",
		b"0000000001111111110011",
		b"0000000010000000001110",
		b"0000000010000000100100",
		b"0000000010000000110101",
		b"0000000010000001000001",
		b"0000000010000001001010",
		b"0000000010000001001101",
		b"0000000010000001001100",
		b"0000000010000001000111",
		b"0000000010000000111101",
		b"0000000010000000101110",
		b"0000000010000000011011",
		b"0000000010000000000100",
		b"0000000001111111101000",
		b"0000000001111111001000",
		b"0000000001111110100011",
		b"0000000001111101111010",
		b"0000000001111101001101",
		b"0000000001111100011011",
		b"0000000001111011100110",
		b"0000000001111010101100",
		b"0000000001111001101110",
		b"0000000001111000101100",
		b"0000000001110111100110",
		b"0000000001110110011100",
		b"0000000001110101001110",
		b"0000000001110011111100",
		b"0000000001110010100111",
		b"0000000001110001001110",
		b"0000000001101111110001",
		b"0000000001101110010000",
		b"0000000001101100101100",
		b"0000000001101011000100",
		b"0000000001101001011001",
		b"0000000001100111101011",
		b"0000000001100101111001",
		b"0000000001100100000100",
		b"0000000001100010001100",
		b"0000000001100000010001",
		b"0000000001011110010011",
		b"0000000001011100010010",
		b"0000000001011010001110",
		b"0000000001011000000111",
		b"0000000001010101111110",
		b"0000000001010011110010",
		b"0000000001010001100100",
		b"0000000001001111010011",
		b"0000000001001101000000",
		b"0000000001001010101011",
		b"0000000001001000010100",
		b"0000000001000101111010",
		b"0000000001000011011111",
		b"0000000001000001000010",
		b"0000000000111110100011",
		b"0000000000111100000010",
		b"0000000000111001011111",
		b"0000000000110110111100",
		b"0000000000110100010110",
		b"0000000000110001110000",
		b"0000000000101111001000",
		b"0000000000101100011111",
		b"0000000000101001110101",
		b"0000000000100111001010",
		b"0000000000100100011110",
		b"0000000000100001110010",
		b"0000000000011111000100",
		b"0000000000011100010111",
		b"0000000000011001101001",
		b"0000000000010110111010",
		b"0000000000010100001011",
		b"0000000000010001011100",
		b"0000000000001110101101",
		b"0000000000001011111110",
		b"0000000000001001001111",
		b"0000000000000110100000",
		b"0000000000000011110010",
		b"0000000000000001000100",
		b"1111111111111110010110",
		b"1111111111111011101010",
		b"1111111111111000111101",
		b"1111111111110110010010",
		b"1111111111110011100111",
		b"1111111111110000111101",
		b"1111111111101110010101",
		b"1111111111101011101101",
		b"1111111111101001000111",
		b"1111111111100110100010",
		b"1111111111100011111110",
		b"1111111111100001011100",
		b"1111111111011110111011",
		b"1111111111011100011100",
		b"1111111111011001111110",
		b"1111111111010111100011",
		b"1111111111010101001001",
		b"1111111111010010110001",
		b"1111111111010000011100",
		b"1111111111001110001000",
		b"1111111111001011110110",
		b"1111111111001001100111",
		b"1111111111000111011010",
		b"1111111111000101010000",
		b"1111111111000011000111",
		b"1111111111000001000010",
		b"1111111110111110111111",
		b"1111111110111100111110",
		b"1111111110111011000000",
		b"1111111110111001000101",
		b"1111111110110111001101",
		b"1111111110110101011000",
		b"1111111110110011100101",
		b"1111111110110001110110",
		b"1111111110110000001001",
		b"1111111110101110100000",
		b"1111111110101100111001",
		b"1111111110101011010110",
		b"1111111110101001110110",
		b"1111111110101000011010",
		b"1111111110100111000000",
		b"1111111110100101101010",
		b"1111111110100100010111",
		b"1111111110100011001000",
		b"1111111110100001111100",
		b"1111111110100000110011",
		b"1111111110011111101110",
		b"1111111110011110101101",
		b"1111111110011101101111",
		b"1111111110011100110100",
		b"1111111110011011111101",
		b"1111111110011011001010",
		b"1111111110011010011010",
		b"1111111110011001101110",
		b"1111111110011001000101",
		b"1111111110011000100000",
		b"1111111110010111111111",
		b"1111111110010111100010",
		b"1111111110010111000111",
		b"1111111110010110110001",
		b"1111111110010110011110",
		b"1111111110010110001111",
		b"1111111110010110000100",
		b"1111111110010101111100",
		b"1111111110010101111000",
		b"1111111110010101110111",
		b"1111111110010101111010",
		b"1111111110010110000001",
		b"1111111110010110001011",
		b"1111111110010110011001",
		b"1111111110010110101010",
		b"1111111110010110111111",
		b"1111111110010111010111",
		b"1111111110010111110011",
		b"1111111110011000010010",
		b"1111111110011000110101",
		b"1111111110011001011011",
		b"1111111110011010000100",
		b"1111111110011010110000",
		b"1111111110011011100000",
		b"1111111110011100010011",
		b"1111111110011101001010",
		b"1111111110011110000011",
		b"1111111110011111000000",
		b"1111111110011111111111",
		b"1111111110100001000010",
		b"1111111110100010001000",
		b"1111111110100011010000",
		b"1111111110100100011100",
		b"1111111110100101101010",
		b"1111111110100110111011",
		b"1111111110101000001111",
		b"1111111110101001100101",
		b"1111111110101010111110",
		b"1111111110101100011010",
		b"1111111110101101111000",
		b"1111111110101111011001",
		b"1111111110110000111100",
		b"1111111110110010100001",
		b"1111111110110100001001",
		b"1111111110110101110010",
		b"1111111110110111011110",
		b"1111111110111001001100",
		b"1111111110111010111100",
		b"1111111110111100101110",
		b"1111111110111110100010",
		b"1111111111000000010111",
		b"1111111111000010001110",
		b"1111111111000100000111",
		b"1111111111000110000010",
		b"1111111111000111111110",
		b"1111111111001001111011",
		b"1111111111001011111010",
		b"1111111111001101111010",
		b"1111111111001111111011",
		b"1111111111010001111101",
		b"1111111111010100000001",
		b"1111111111010110000101",
		b"1111111111011000001011",
		b"1111111111011010010001",
		b"1111111111011100011000",
		b"1111111111011110011111",
		b"1111111111100000101000",
		b"1111111111100010110001",
		b"1111111111100100111010",
		b"1111111111100111000100",
		b"1111111111101001001110",
		b"1111111111101011011000",
		b"1111111111101101100010",
		b"1111111111101111101101",
		b"1111111111110001110111",
		b"1111111111110100000001",
		b"1111111111110110001100",
		b"1111111111111000010110",
		b"1111111111111010100000",
		b"1111111111111100101001",
		b"1111111111111110110010",
		b"0000000000000000111011",
		b"0000000000000011000010",
		b"0000000000000101001010",
		b"0000000000000111010000",
		b"0000000000001001010110",
		b"0000000000001011011011",
		b"0000000000001101011111",
		b"0000000000001111100010",
		b"0000000000010001100100",
		b"0000000000010011100100",
		b"0000000000010101100100",
		b"0000000000010111100010",
		b"0000000000011001011111",
		b"0000000000011011011011",
		b"0000000000011101010101",
		b"0000000000011111001110",
		b"0000000000100001000101",
		b"0000000000100010111010",
		b"0000000000100100101110",
		b"0000000000100110100000",
		b"0000000000101000010000",
		b"0000000000101001111111",
		b"0000000000101011101011",
		b"0000000000101101010110",
		b"0000000000101110111110",
		b"0000000000110000100101",
		b"0000000000110010001001",
		b"0000000000110011101011",
		b"0000000000110101001011",
		b"0000000000110110101001",
		b"0000000000111000000101",
		b"0000000000111001011110",
		b"0000000000111010110101",
		b"0000000000111100001001",
		b"0000000000111101011011",
		b"0000000000111110101010",
		b"0000000000111111110111",
		b"0000000001000001000010",
		b"0000000001000010001010",
		b"0000000001000011001111",
		b"0000000001000100010001",
		b"0000000001000101010001",
		b"0000000001000110001110",
		b"0000000001000111001001",
		b"0000000001001000000001",
		b"0000000001001000110110",
		b"0000000001001001101000",
		b"0000000001001010011000",
		b"0000000001001011000100",
		b"0000000001001011101110",
		b"0000000001001100010101",
		b"0000000001001100111001",
		b"0000000001001101011010",
		b"0000000001001101111001",
		b"0000000001001110010100",
		b"0000000001001110101101",
		b"0000000001001111000011",
		b"0000000001001111010110",
		b"0000000001001111100110",
		b"0000000001001111110011",
		b"0000000001001111111101",
		b"0000000001010000000101",
		b"0000000001010000001001",
		b"0000000001010000001011",
		b"0000000001010000001010",
		b"0000000001010000000110",
		b"0000000001001111111111",
		b"0000000001001111110101",
		b"0000000001001111101001",
		b"0000000001001111011010",
		b"0000000001001111001000",
		b"0000000001001110110011",
		b"0000000001001110011011",
		b"0000000001001110000001",
		b"0000000001001101100100",
		b"0000000001001101000101",
		b"0000000001001100100010",
		b"0000000001001011111110",
		b"0000000001001011010110",
		b"0000000001001010101100",
		b"0000000001001010000000",
		b"0000000001001001010001",
		b"0000000001001000011111",
		b"0000000001000111101100",
		b"0000000001000110110101",
		b"0000000001000101111101",
		b"0000000001000101000010",
		b"0000000001000100000101",
		b"0000000001000011000101",
		b"0000000001000010000100",
		b"0000000001000001000000",
		b"0000000000111111111010",
		b"0000000000111110110011",
		b"0000000000111101101001",
		b"0000000000111100011101",
		b"0000000000111011001111",
		b"0000000000111001111111",
		b"0000000000111000101110",
		b"0000000000110111011011",
		b"0000000000110110000110",
		b"0000000000110100101111",
		b"0000000000110011010111",
		b"0000000000110001111101",
		b"0000000000110000100010",
		b"0000000000101111000101",
		b"0000000000101101100111",
		b"0000000000101100000111",
		b"0000000000101010100110",
		b"0000000000101001000100",
		b"0000000000100111100001",
		b"0000000000100101111101",
		b"0000000000100100010111",
		b"0000000000100010110001",
		b"0000000000100001001001",
		b"0000000000011111100001",
		b"0000000000011101110111",
		b"0000000000011100001110",
		b"0000000000011010100011",
		b"0000000000011000110111",
		b"0000000000010111001011",
		b"0000000000010101011111",
		b"0000000000010011110010",
		b"0000000000010010000100",
		b"0000000000010000010111",
		b"0000000000001110101001",
		b"0000000000001100111010",
		b"0000000000001011001100",
		b"0000000000001001011101",
		b"0000000000000111101110",
		b"0000000000000101111111",
		b"0000000000000100010001",
		b"0000000000000010100010",
		b"0000000000000000110100",
		b"1111111111111111000101",
		b"1111111111111101010111",
		b"1111111111111011101010",
		b"1111111111111001111101",
		b"1111111111111000010000",
		b"1111111111110110100100",
		b"1111111111110100111000",
		b"1111111111110011001101",
		b"1111111111110001100010",
		b"1111111111101111111001",
		b"1111111111101110010000",
		b"1111111111101100101000",
		b"1111111111101011000000",
		b"1111111111101001011010",
		b"1111111111100111110101",
		b"1111111111100110010000",
		b"1111111111100100101101",
		b"1111111111100011001011",
		b"1111111111100001101010",
		b"1111111111100000001011",
		b"1111111111011110101100",
		b"1111111111011101001111",
		b"1111111111011011110011",
		b"1111111111011010011001",
		b"1111111111011001000000",
		b"1111111111010111101001",
		b"1111111111010110010011",
		b"1111111111010100111111",
		b"1111111111010011101100",
		b"1111111111010010011011",
		b"1111111111010001001100",
		b"1111111111001111111110",
		b"1111111111001110110010",
		b"1111111111001101101000",
		b"1111111111001100100000",
		b"1111111111001011011010",
		b"1111111111001010010101",
		b"1111111111001001010011",
		b"1111111111001000010010",
		b"1111111111000111010011",
		b"1111111111000110010111",
		b"1111111111000101011100",
		b"1111111111000100100011",
		b"1111111111000011101101",
		b"1111111111000010111000",
		b"1111111111000010000110",
		b"1111111111000001010110",
		b"1111111111000000101000",
		b"1111111110111111111100",
		b"1111111110111111010010",
		b"1111111110111110101010",
		b"1111111110111110000101",
		b"1111111110111101100010",
		b"1111111110111101000001",
		b"1111111110111100100010",
		b"1111111110111100000110",
		b"1111111110111011101100",
		b"1111111110111011010100",
		b"1111111110111010111110",
		b"1111111110111010101011",
		b"1111111110111010011001",
		b"1111111110111010001011",
		b"1111111110111001111110",
		b"1111111110111001110100",
		b"1111111110111001101011",
		b"1111111110111001100110",
		b"1111111110111001100010",
		b"1111111110111001100001",
		b"1111111110111001100010",
		b"1111111110111001100101",
		b"1111111110111001101010",
		b"1111111110111001110010",
		b"1111111110111001111011",
		b"1111111110111010000111",
		b"1111111110111010010101",
		b"1111111110111010100110",
		b"1111111110111010111000",
		b"1111111110111011001100",
		b"1111111110111011100011",
		b"1111111110111011111100",
		b"1111111110111100010110",
		b"1111111110111100110011",
		b"1111111110111101010010",
		b"1111111110111101110011",
		b"1111111110111110010110",
		b"1111111110111110111010",
		b"1111111110111111100001",
		b"1111111111000000001001",
		b"1111111111000000110100",
		b"1111111111000001100000",
		b"1111111111000010001110",
		b"1111111111000010111110",
		b"1111111111000011101111",
		b"1111111111000100100010",
		b"1111111111000101010111",
		b"1111111111000110001110",
		b"1111111111000111000110",
		b"1111111111001000000000",
		b"1111111111001000111011",
		b"1111111111001001110111",
		b"1111111111001010110110",
		b"1111111111001011110101",
		b"1111111111001100110110",
		b"1111111111001101111000",
		b"1111111111001110111100",
		b"1111111111010000000001",
		b"1111111111010001000111",
		b"1111111111010010001110",
		b"1111111111010011010110",
		b"1111111111010100100000",
		b"1111111111010101101010",
		b"1111111111010110110110",
		b"1111111111011000000010",
		b"1111111111011001010000",
		b"1111111111011010011110",
		b"1111111111011011101101",
		b"1111111111011100111101",
		b"1111111111011110001110",
		b"1111111111011111011111",
		b"1111111111100000110001",
		b"1111111111100010000011",
		b"1111111111100011010110",
		b"1111111111100100101010",
		b"1111111111100101111110",
		b"1111111111100111010011",
		b"1111111111101000100111",
		b"1111111111101001111101",
		b"1111111111101011010010",
		b"1111111111101100101000",
		b"1111111111101101111110",
		b"1111111111101111010100",
		b"1111111111110000101010",
		b"1111111111110010000000",
		b"1111111111110011010110",
		b"1111111111110100101100",
		b"1111111111110110000010",
		b"1111111111110111011000",
		b"1111111111111000101101",
		b"1111111111111010000011",
		b"1111111111111011011000",
		b"1111111111111100101101",
		b"1111111111111110000001",
		b"1111111111111111010101",
		b"0000000000000000101001",
		b"0000000000000001111100",
		b"0000000000000011001111",
		b"0000000000000100100001",
		b"0000000000000101110010",
		b"0000000000000111000011",
		b"0000000000001000010011",
		b"0000000000001001100010",
		b"0000000000001010110001",
		b"0000000000001011111110",
		b"0000000000001101001011",
		b"0000000000001110010111",
		b"0000000000001111100010",
		b"0000000000010000101100",
		b"0000000000010001110101",
		b"0000000000010010111101",
		b"0000000000010100000100",
		b"0000000000010101001010",
		b"0000000000010110001111",
		b"0000000000010111010010",
		b"0000000000011000010100",
		b"0000000000011001010101",
		b"0000000000011010010101",
		b"0000000000011011010011",
		b"0000000000011100010001",
		b"0000000000011101001100",
		b"0000000000011110000111",
		b"0000000000011111000000",
		b"0000000000011111110111",
		b"0000000000100000101101",
		b"0000000000100001100010",
		b"0000000000100010010101",
		b"0000000000100011000110",
		b"0000000000100011110110",
		b"0000000000100100100101",
		b"0000000000100101010001",
		b"0000000000100101111101",
		b"0000000000100110100110",
		b"0000000000100111001110",
		b"0000000000100111110100",
		b"0000000000101000011001",
		b"0000000000101000111100",
		b"0000000000101001011101",
		b"0000000000101001111100",
		b"0000000000101010011010",
		b"0000000000101010110110",
		b"0000000000101011010000",
		b"0000000000101011101000",
		b"0000000000101011111111",
		b"0000000000101100010100",
		b"0000000000101100100111",
		b"0000000000101100111000",
		b"0000000000101101001000",
		b"0000000000101101010101",
		b"0000000000101101100001",
		b"0000000000101101101011",
		b"0000000000101101110100",
		b"0000000000101101111010",
		b"0000000000101101111111",
		b"0000000000101110000010",
		b"0000000000101110000011",
		b"0000000000101110000010",
		b"0000000000101110000000",
		b"0000000000101101111100",
		b"0000000000101101110110",
		b"0000000000101101101110",
		b"0000000000101101100101",
		b"0000000000101101011001",
		b"0000000000101101001101",
		b"0000000000101100111110",
		b"0000000000101100101110",
		b"0000000000101100011100",
		b"0000000000101100001000",
		b"0000000000101011110010",
		b"0000000000101011011011",
		b"0000000000101011000011",
		b"0000000000101010101000",
		b"0000000000101010001101",
		b"0000000000101001101111",
		b"0000000000101001010000",
		b"0000000000101000110000",
		b"0000000000101000001101",
		b"0000000000100111101010",
		b"0000000000100111000101",
		b"0000000000100110011110",
		b"0000000000100101110110",
		b"0000000000100101001101",
		b"0000000000100100100010",
		b"0000000000100011110110",
		b"0000000000100011001001",
		b"0000000000100010011010",
		b"0000000000100001101010",
		b"0000000000100000111001",
		b"0000000000100000000111",
		b"0000000000011111010011",
		b"0000000000011110011110",
		b"0000000000011101101000",
		b"0000000000011100110001",
		b"0000000000011011111001",
		b"0000000000011011000000",
		b"0000000000011010000110",
		b"0000000000011001001011",
		b"0000000000011000001111",
		b"0000000000010111010010",
		b"0000000000010110010101",
		b"0000000000010101010110",
		b"0000000000010100010111",
		b"0000000000010011010110",
		b"0000000000010010010101",
		b"0000000000010001010100",
		b"0000000000010000010010",
		b"0000000000001111001111",
		b"0000000000001110001011",
		b"0000000000001101000111",
		b"0000000000001100000010",
		b"0000000000001010111101",
		b"0000000000001001111000",
		b"0000000000001000110010",
		b"0000000000000111101011",
		b"0000000000000110100101",
		b"0000000000000101011110",
		b"0000000000000100010111",
		b"0000000000000011001111",
		b"0000000000000010000111",
		b"0000000000000001000000",
		b"1111111111111111111000",
		b"1111111111111110101111",
		b"1111111111111101100111",
		b"1111111111111100011111",
		b"1111111111111011010111",
		b"1111111111111010001111",
		b"1111111111111001000111",
		b"1111111111110111111111",
		b"1111111111110110111000",
		b"1111111111110101110000",
		b"1111111111110100101001",
		b"1111111111110011100010",
		b"1111111111110010011011",
		b"1111111111110001010101",
		b"1111111111110000001111",
		b"1111111111101111001001",
		b"1111111111101110000100",
		b"1111111111101100111111",
		b"1111111111101011111011",
		b"1111111111101010111000",
		b"1111111111101001110101",
		b"1111111111101000110010",
		b"1111111111100111110000",
		b"1111111111100110101111",
		b"1111111111100101101111",
		b"1111111111100100101111",
		b"1111111111100011110000",
		b"1111111111100010110010",
		b"1111111111100001110100",
		b"1111111111100000111000",
		b"1111111111011111111100",
		b"1111111111011111000001",
		b"1111111111011110000111",
		b"1111111111011101001110",
		b"1111111111011100010110",
		b"1111111111011011011111",
		b"1111111111011010101001",
		b"1111111111011001110100",
		b"1111111111011001000000",
		b"1111111111011000001101",
		b"1111111111010111011011",
		b"1111111111010110101011",
		b"1111111111010101111011",
		b"1111111111010101001101",
		b"1111111111010100100000",
		b"1111111111010011110100",
		b"1111111111010011001001",
		b"1111111111010010100000",
		b"1111111111010001111000",
		b"1111111111010001010001",
		b"1111111111010000101011",
		b"1111111111010000000111",
		b"1111111111001111100100",
		b"1111111111001111000010",
		b"1111111111001110100001",
		b"1111111111001110000010",
		b"1111111111001101100101",
		b"1111111111001101001000",
		b"1111111111001100101110",
		b"1111111111001100010100",
		b"1111111111001011111100",
		b"1111111111001011100101",
		b"1111111111001011010000",
		b"1111111111001010111100",
		b"1111111111001010101001",
		b"1111111111001010011000",
		b"1111111111001010001001",
		b"1111111111001001111011",
		b"1111111111001001101110",
		b"1111111111001001100010",
		b"1111111111001001011001",
		b"1111111111001001010000",
		b"1111111111001001001001",
		b"1111111111001001000011",
		b"1111111111001000111111",
		b"1111111111001000111101",
		b"1111111111001000111011",
		b"1111111111001000111011",
		b"1111111111001000111101",
		b"1111111111001001000000",
		b"1111111111001001000100",
		b"1111111111001001001010",
		b"1111111111001001010001",
		b"1111111111001001011001",
		b"1111111111001001100011",
		b"1111111111001001101111",
		b"1111111111001001111011",
		b"1111111111001010001001",
		b"1111111111001010011000",
		b"1111111111001010101001",
		b"1111111111001010111011",
		b"1111111111001011001110",
		b"1111111111001011100010",
		b"1111111111001011111000",
		b"1111111111001100001111",
		b"1111111111001100100111",
		b"1111111111001101000000",
		b"1111111111001101011011",
		b"1111111111001101110111",
		b"1111111111001110010100",
		b"1111111111001110110010",
		b"1111111111001111010001",
		b"1111111111001111110001",
		b"1111111111010000010011",
		b"1111111111010000110101",
		b"1111111111010001011000",
		b"1111111111010001111101",
		b"1111111111010010100010",
		b"1111111111010011001001",
		b"1111111111010011110000",
		b"1111111111010100011001",
		b"1111111111010101000010",
		b"1111111111010101101100",
		b"1111111111010110010111",
		b"1111111111010111000011",
		b"1111111111010111110000",
		b"1111111111011000011101",
		b"1111111111011001001011",
		b"1111111111011001111010",
		b"1111111111011010101010",
		b"1111111111011011011010",
		b"1111111111011100001011",
		b"1111111111011100111101",
		b"1111111111011101101111",
		b"1111111111011110100010",
		b"1111111111011111010101",
		b"1111111111100000001001",
		b"1111111111100000111101",
		b"1111111111100001110010",
		b"1111111111100010100111",
		b"1111111111100011011101",
		b"1111111111100100010011",
		b"1111111111100101001001",
		b"1111111111100110000000",
		b"1111111111100110110111",
		b"1111111111100111101110",
		b"1111111111101000100110",
		b"1111111111101001011101",
		b"1111111111101010010101",
		b"1111111111101011001101",
		b"1111111111101100000101",
		b"1111111111101100111101",
		b"1111111111101101110110",
		b"1111111111101110101110",
		b"1111111111101111100110",
		b"1111111111110000011111",
		b"1111111111110001010111",
		b"1111111111110010001111",
		b"1111111111110011000111",
		b"1111111111110011111111",
		b"1111111111110100110111",
		b"1111111111110101101110",
		b"1111111111110110100101",
		b"1111111111110111011100",
		b"1111111111111000010011",
		b"1111111111111001001010",
		b"1111111111111010000000",
		b"1111111111111010110110",
		b"1111111111111011101011",
		b"1111111111111100100000",
		b"1111111111111101010100",
		b"1111111111111110001000",
		b"1111111111111110111100",
		b"1111111111111111101111",
		b"0000000000000000100010",
		b"0000000000000001010100",
		b"0000000000000010000101",
		b"0000000000000010110110",
		b"0000000000000011100110",
		b"0000000000000100010101",
		b"0000000000000101000100",
		b"0000000000000101110010",
		b"0000000000000110011111",
		b"0000000000000111001100",
		b"0000000000000111111000",
		b"0000000000001000100011",
		b"0000000000001001001101",
		b"0000000000001001110111",
		b"0000000000001010011111",
		b"0000000000001011000111",
		b"0000000000001011101110",
		b"0000000000001100010011",
		b"0000000000001100111000",
		b"0000000000001101011100",
		b"0000000000001110000000",
		b"0000000000001110100010",
		b"0000000000001111000011",
		b"0000000000001111100011",
		b"0000000000010000000010",
		b"0000000000010000100000",
		b"0000000000010000111101",
		b"0000000000010001011001",
		b"0000000000010001110100",
		b"0000000000010010001101",
		b"0000000000010010100110",
		b"0000000000010010111110",
		b"0000000000010011010100",
		b"0000000000010011101010",
		b"0000000000010011111110",
		b"0000000000010100010001",
		b"0000000000010100100011",
		b"0000000000010100110011",
		b"0000000000010101000011",
		b"0000000000010101010001",
		b"0000000000010101011110",
		b"0000000000010101101010",
		b"0000000000010101110101",
		b"0000000000010101111111",
		b"0000000000010110000111",
		b"0000000000010110001110",
		b"0000000000010110010100",
		b"0000000000010110011001",
		b"0000000000010110011101",
		b"0000000000010110011111",
		b"0000000000010110100000",
		b"0000000000010110100000",
		b"0000000000010110011110",
		b"0000000000010110011100",
		b"0000000000010110011000",
		b"0000000000010110010011",
		b"0000000000010110001101",
		b"0000000000010110000110",
		b"0000000000010101111101",
		b"0000000000010101110011",
		b"0000000000010101101000",
		b"0000000000010101011100",
		b"0000000000010101001111",
		b"0000000000010101000000",
		b"0000000000010100110000",
		b"0000000000010100011111",
		b"0000000000010100001101",
		b"0000000000010011111010",
		b"0000000000010011100110",
		b"0000000000010011010000",
		b"0000000000010010111010",
		b"0000000000010010100010",
		b"0000000000010010001001",
		b"0000000000010001101111",
		b"0000000000010001010100",
		b"0000000000010000111000",
		b"0000000000010000011011",
		b"0000000000001111111101",
		b"0000000000001111011110",
		b"0000000000001110111101",
		b"0000000000001110011100",
		b"0000000000001101111010",
		b"0000000000001101010111",
		b"0000000000001100110011",
		b"0000000000001100001110",
		b"0000000000001011101000",
		b"0000000000001011000001",
		b"0000000000001010011001",
		b"0000000000001001110000",
		b"0000000000001001000111",
		b"0000000000001000011100",
		b"0000000000000111110001",
		b"0000000000000111000101",
		b"0000000000000110011000",
		b"0000000000000101101011",
		b"0000000000000100111100",
		b"0000000000000100001101",
		b"0000000000000011011101",
		b"0000000000000010101101",
		b"0000000000000001111100",
		b"0000000000000001001010",
		b"0000000000000000011000",
		b"1111111111111111100101",
		b"1111111111111110110001",
		b"1111111111111101111101",
		b"1111111111111101001000",
		b"1111111111111100010011",
		b"1111111111111011011101",
		b"1111111111111010100111",
		b"1111111111111001110000",
		b"1111111111111000111001",
		b"1111111111111000000001",
		b"1111111111110111001001",
		b"1111111111110110010001",
		b"1111111111110101011000",
		b"1111111111110100011111",
		b"1111111111110011100110",
		b"1111111111110010101100",
		b"1111111111110001110010",
		b"1111111111110000111000",
		b"1111111111101111111110",
		b"1111111111101111000011",
		b"1111111111101110001001",
		b"1111111111101101001110",
		b"1111111111101100010011",
		b"1111111111101011011000",
		b"1111111111101010011101",
		b"1111111111101001100001",
		b"1111111111101000100110",
		b"1111111111100111101011",
		b"1111111111100110110000",
		b"1111111111100101110100",
		b"1111111111100100111001",
		b"1111111111100011111110",
		b"1111111111100011000011",
		b"1111111111100010001000",
		b"1111111111100001001110",
		b"1111111111100000010011",
		b"1111111111011111011001",
		b"1111111111011110011111",
		b"1111111111011101100101",
		b"1111111111011100101011",
		b"1111111111011011110010",
		b"1111111111011010111001",
		b"1111111111011010000000",
		b"1111111111011001001000",
		b"1111111111011000010000",
		b"1111111111010111011000",
		b"1111111111010110100001",
		b"1111111111010101101010",
		b"1111111111010100110100",
		b"1111111111010011111110",
		b"1111111111010011001000",
		b"1111111111010010010100",
		b"1111111111010001011111",
		b"1111111111010000101011",
		b"1111111111001111111000",
		b"1111111111001111000101",
		b"1111111111001110010011",
		b"1111111111001101100001",
		b"1111111111001100110000",
		b"1111111111001100000000",
		b"1111111111001011010000",
		b"1111111111001010100001",
		b"1111111111001001110011",
		b"1111111111001001000110",
		b"1111111111001000011001",
		b"1111111111000111101100",
		b"1111111111000111000001",
		b"1111111111000110010110",
		b"1111111111000101101101",
		b"1111111111000101000100",
		b"1111111111000100011011",
		b"1111111111000011110100",
		b"1111111111000011001101",
		b"1111111111000010100111",
		b"1111111111000010000010",
		b"1111111111000001011110",
		b"1111111111000000111011",
		b"1111111111000000011001",
		b"1111111110111111110111",
		b"1111111110111111010111",
		b"1111111110111110110111",
		b"1111111110111110011001",
		b"1111111110111101111011",
		b"1111111110111101011110",
		b"1111111110111101000010",
		b"1111111110111100100111",
		b"1111111110111100001110",
		b"1111111110111011110101",
		b"1111111110111011011101",
		b"1111111110111011000110",
		b"1111111110111010110000",
		b"1111111110111010011011",
		b"1111111110111010000111",
		b"1111111110111001110100",
		b"1111111110111001100010",
		b"1111111110111001010001",
		b"1111111110111001000001",
		b"1111111110111000110010",
		b"1111111110111000100100",
		b"1111111110111000010111",
		b"1111111110111000001011",
		b"1111111110111000000001",
		b"1111111110110111110111",
		b"1111111110110111101110",
		b"1111111110110111100110",
		b"1111111110110111100000",
		b"1111111110110111011010",
		b"1111111110110111010101",
		b"1111111110110111010010",
		b"1111111110110111001111",
		b"1111111110110111001110",
		b"1111111110110111001101",
		b"1111111110110111001110",
		b"1111111110110111001111",
		b"1111111110110111010010",
		b"1111111110110111010101",
		b"1111111110110111011010",
		b"1111111110110111100000",
		b"1111111110110111100110",
		b"1111111110110111101110",
		b"1111111110110111110110",
		b"1111111110111000000000",
		b"1111111110111000001011",
		b"1111111110111000010110",
		b"1111111110111000100011",
		b"1111111110111000110000",
		b"1111111110111000111110",
		b"1111111110111001001110",
		b"1111111110111001011110",
		b"1111111110111001101111",
		b"1111111110111010000010",
		b"1111111110111010010101",
		b"1111111110111010101001",
		b"1111111110111010111110",
		b"1111111110111011010100",
		b"1111111110111011101010",
		b"1111111110111100000010",
		b"1111111110111100011010",
		b"1111111110111100110011",
		b"1111111110111101001110",
		b"1111111110111101101001",
		b"1111111110111110000100",
		b"1111111110111110100001",
		b"1111111110111110111110",
		b"1111111110111111011100",
		b"1111111110111111111011",
		b"1111111111000000011011",
		b"1111111111000000111100",
		b"1111111111000001011101",
		b"1111111111000001111111",
		b"1111111111000010100001",
		b"1111111111000011000101",
		b"1111111111000011101001",
		b"1111111111000100001110",
		b"1111111111000100110011",
		b"1111111111000101011001",
		b"1111111111000110000000",
		b"1111111111000110100111",
		b"1111111111000111001111",
		b"1111111111000111110111",
		b"1111111111001000100000",
		b"1111111111001001001010",
		b"1111111111001001110100",
		b"1111111111001010011111",
		b"1111111111001011001010",
		b"1111111111001011110110",
		b"1111111111001100100010",
		b"1111111111001101001111",
		b"1111111111001101111100",
		b"1111111111001110101010",
		b"1111111111001111011000",
		b"1111111111010000000111",
		b"1111111111010000110110",
		b"1111111111010001100101",
		b"1111111111010010010101",
		b"1111111111010011000101",
		b"1111111111010011110101",
		b"1111111111010100100110",
		b"1111111111010101010111",
		b"1111111111010110001000",
		b"1111111111010110111010",
		b"1111111111010111101100",
		b"1111111111011000011110",
		b"1111111111011001010000",
		b"1111111111011010000011",
		b"1111111111011010110110",
		b"1111111111011011101001",
		b"1111111111011100011100",
		b"1111111111011101010000",
		b"1111111111011110000011",
		b"1111111111011110110111",
		b"1111111111011111101011",
		b"1111111111100000011111",
		b"1111111111100001010011",
		b"1111111111100010000111",
		b"1111111111100010111011",
		b"1111111111100011110000",
		b"1111111111100100100100",
		b"1111111111100101011000",
		b"1111111111100110001101",
		b"1111111111100111000001",
		b"1111111111100111110101",
		b"1111111111101000101010",
		b"1111111111101001011110",
		b"1111111111101010010010",
		b"1111111111101011000110",
		b"1111111111101011111010",
		b"1111111111101100101110",
		b"1111111111101101100010",
		b"1111111111101110010110",
		b"1111111111101111001001",
		b"1111111111101111111101",
		b"1111111111110000110000",
		b"1111111111110001100011",
		b"1111111111110010010110",
		b"1111111111110011001001",
		b"1111111111110011111011",
		b"1111111111110100101101",
		b"1111111111110101100000",
		b"1111111111110110010001",
		b"1111111111110111000011",
		b"1111111111110111110100",
		b"1111111111111000100101",
		b"1111111111111001010110",
		b"1111111111111010000110",
		b"1111111111111010110111",
		b"1111111111111011100110",
		b"1111111111111100010110",
		b"1111111111111101000101",
		b"1111111111111101110100",
		b"1111111111111110100010",
		b"1111111111111111010001",
		b"1111111111111111111110",
		b"0000000000000000101100",
		b"0000000000000001011001",
		b"0000000000000010000101",
		b"0000000000000010110001",
		b"0000000000000011011101",
		b"0000000000000100001001",
		b"0000000000000100110100",
		b"0000000000000101011110",
		b"0000000000000110001000",
		b"0000000000000110110010",
		b"0000000000000111011011",
		b"0000000000001000000011",
		b"0000000000001000101100",
		b"0000000000001001010011",
		b"0000000000001001111011",
		b"0000000000001010100001",
		b"0000000000001011001000",
		b"0000000000001011101101",
		b"0000000000001100010011",
		b"0000000000001100111000",
		b"0000000000001101011100",
		b"0000000000001110000000",
		b"0000000000001110100011",
		b"0000000000001111000110",
		b"0000000000001111101000",
		b"0000000000010000001001",
		b"0000000000010000101010",
		b"0000000000010001001011",
		b"0000000000010001101011",
		b"0000000000010010001011",
		b"0000000000010010101001",
		b"0000000000010011001000",
		b"0000000000010011100110",
		b"0000000000010100000011",
		b"0000000000010100100000",
		b"0000000000010100111100",
		b"0000000000010101011000",
		b"0000000000010101110011",
		b"0000000000010110001101",
		b"0000000000010110100111",
		b"0000000000010111000000",
		b"0000000000010111011001",
		b"0000000000010111110010",
		b"0000000000011000001001",
		b"0000000000011000100000",
		b"0000000000011000110111",
		b"0000000000011001001101",
		b"0000000000011001100010",
		b"0000000000011001110111",
		b"0000000000011010001100",
		b"0000000000011010011111",
		b"0000000000011010110010",
		b"0000000000011011000101",
		b"0000000000011011010111",
		b"0000000000011011101001",
		b"0000000000011011111010",
		b"0000000000011100001010",
		b"0000000000011100011010",
		b"0000000000011100101001",
		b"0000000000011100111000",
		b"0000000000011101000110",
		b"0000000000011101010100",
		b"0000000000011101100001",
		b"0000000000011101101110",
		b"0000000000011101111010",
		b"0000000000011110000110",
		b"0000000000011110010001",
		b"0000000000011110011011",
		b"0000000000011110100101",
		b"0000000000011110101111",
		b"0000000000011110111000",
		b"0000000000011111000000",
		b"0000000000011111001000",
		b"0000000000011111010000",
		b"0000000000011111010111",
		b"0000000000011111011101",
		b"0000000000011111100011",
		b"0000000000011111101001",
		b"0000000000011111101110",
		b"0000000000011111110010",
		b"0000000000011111110110",
		b"0000000000011111111010",
		b"0000000000011111111101",
		b"0000000000100000000000",
		b"0000000000100000000010",
		b"0000000000100000000100",
		b"0000000000100000000110",
		b"0000000000100000000111",
		b"0000000000100000000111",
		b"0000000000100000000111",
		b"0000000000100000000111",
		b"0000000000100000000110",
		b"0000000000100000000101",
		b"0000000000100000000100",
		b"0000000000100000000010",
		b"0000000000100000000000",
		b"0000000000011111111101",
		b"0000000000011111111010",
		b"0000000000011111110111",
		b"0000000000011111110011",
		b"0000000000011111101111",
		b"0000000000011111101010",
		b"0000000000011111100110",
		b"0000000000011111100000",
		b"0000000000011111011011",
		b"0000000000011111010101",
		b"0000000000011111001111",
		b"0000000000011111001001",
		b"0000000000011111000010",
		b"0000000000011110111011",
		b"0000000000011110110011",
		b"0000000000011110101100",
		b"0000000000011110100100",
		b"0000000000011110011100",
		b"0000000000011110010011",
		b"0000000000011110001010",
		b"0000000000011110000001",
		b"0000000000011101111000",
		b"0000000000011101101111",
		b"0000000000011101100101",
		b"0000000000011101011011",
		b"0000000000011101010001",
		b"0000000000011101000110",
		b"0000000000011100111100",
		b"0000000000011100110001",
		b"0000000000011100100110",
		b"0000000000011100011011",
		b"0000000000011100001111",
		b"0000000000011100000011",
		b"0000000000011011111000",
		b"0000000000011011101100",
		b"0000000000011011011111",
		b"0000000000011011010011",
		b"0000000000011011000111",
		b"0000000000011010111010",
		b"0000000000011010101101",
		b"0000000000011010100000",
		b"0000000000011010010011",
		b"0000000000011010000110",
		b"0000000000011001111001",
		b"0000000000011001101011",
		b"0000000000011001011110",
		b"0000000000011001010000",
		b"0000000000011001000010",
		b"0000000000011000110100",
		b"0000000000011000100110",
		b"0000000000011000011000",
		b"0000000000011000001010",
		b"0000000000010111111100",
		b"0000000000010111101110",
		b"0000000000010111011111",
		b"0000000000010111010001",
		b"0000000000010111000011",
		b"0000000000010110110100",
		b"0000000000010110100110",
		b"0000000000010110010111",
		b"0000000000010110001000",
		b"0000000000010101111010",
		b"0000000000010101101011",
		b"0000000000010101011100",
		b"0000000000010101001101",
		b"0000000000010100111111",
		b"0000000000010100110000",
		b"0000000000010100100001",
		b"0000000000010100010010",
		b"0000000000010100000100",
		b"0000000000010011110101",
		b"0000000000010011100110",
		b"0000000000010011010111",
		b"0000000000010011001001",
		b"0000000000010010111010",
		b"0000000000010010101011",
		b"0000000000010010011100",
		b"0000000000010010001110",
		b"0000000000010001111111",
		b"0000000000010001110001",
		b"0000000000010001100010",
		b"0000000000010001010100",
		b"0000000000010001000101",
		b"0000000000010000110111",
		b"0000000000010000101000",
		b"0000000000010000011010",
		b"0000000000010000001100",
		b"0000000000001111111110",
		b"0000000000001111110000",
		b"0000000000001111100010",
		b"0000000000001111010100",
		b"0000000000001111000110",
		b"0000000000001110111000",
		b"0000000000001110101010",
		b"0000000000001110011100",
		b"0000000000001110001111",
		b"0000000000001110000001",
		b"0000000000001101110100",
		b"0000000000001101100111",
		b"0000000000001101011001",
		b"0000000000001101001100",
		b"0000000000001100111111",
		b"0000000000001100110010",
		b"0000000000001100100101",
		b"0000000000001100011001",
		b"0000000000001100001100",
		b"0000000000001011111111",
		b"0000000000001011110011",
		b"0000000000001011100110",
		b"0000000000001011011010",
		b"0000000000001011001110",
		b"0000000000001011000010",
		b"0000000000001010110110",
		b"0000000000001010101010",
		b"0000000000001010011111",
		b"0000000000001010010011",
		b"0000000000001010000111",
		b"0000000000001001111100",
		b"0000000000001001110001",
		b"0000000000001001100110",
		b"0000000000001001011011",
		b"0000000000001001010000",
		b"0000000000001001000101",
		b"0000000000001000111010",
		b"0000000000001000110000",
		b"0000000000001000100101",
		b"0000000000001000011011",
		b"0000000000001000010001",
		b"0000000000001000000111",
		b"0000000000000111111101",
		b"0000000000000111110011",
		b"0000000000000111101001",
		b"0000000000000111100000",
		b"0000000000000111010110",
		b"0000000000000111001101",
		b"0000000000000111000011",
		b"0000000000000110111010",
		b"0000000000000110110001",
		b"0000000000000110101000",
		b"0000000000000110100000",
		b"0000000000000110010111",
		b"0000000000000110001111",
		b"0000000000000110000110",
		b"0000000000000101111110",
		b"0000000000000101110110",
		b"0000000000000101101110",
		b"0000000000000101100110",
		b"0000000000000101011110",
		b"0000000000000101010110",
		b"0000000000000101001111",
		b"0000000000000101000111",
		b"0000000000000101000000",
		b"0000000000000100111001",
		b"0000000000000100110010",
		b"0000000000000100101011",
		b"0000000000000100100100",
		b"0000000000000100011101",
		b"0000000000000100010110",
		b"0000000000000100010000",
		b"0000000000000100001001",
		b"0000000000000100000011",
		b"0000000000000011111101",
		b"0000000000000011110111",
		b"0000000000000011110001",
		b"0000000000000011101011",
		b"0000000000000011100101",
		b"0000000000000011011111",
		b"0000000000000011011010",
		b"0000000000000011010100",
		b"0000000000000011001111",
		b"0000000000000011001010",
		b"0000000000000011000100",
		b"0000000000000010111111",
		b"0000000000000010111010",
		b"0000000000000010110101",
		b"0000000000000010110001",
		b"0000000000000010101100",
		b"0000000000000010100111",
		b"0000000000000010100011",
		b"0000000000000010011110",
		b"0000000000000010011010",
		b"0000000000000010010110",
		b"0000000000000010010010",
		b"0000000000000010001110",
		b"0000000000000010001010",
		b"0000000000000010000110",
		b"0000000000000010000010",
		b"0000000000000001111110",
		b"0000000000000001111011",
		b"0000000000000001110111",
		b"0000000000000001110011",
		b"0000000000000001110000",
		b"0000000000000001101101",
		b"0000000000000001101001",
		b"0000000000000001100110",
		b"0000000000000001100011",
		b"0000000000000001100000",
		b"0000000000000001011101",
		b"0000000000000001011010",
		b"0000000000000001010111",
		b"0000000000000001010101",
		b"0000000000000001010010",
		b"0000000000000001001111",
		b"0000000000000001001101",
		b"0000000000000001001010",
		b"0000000000000001001000",
		b"0000000000000001000110",
		b"0000000000000001000011",
		b"0000000000000001000001",
		b"0000000000000000111111",
		b"0000000000000000111101",
		b"0000000000000000111011",
		b"0000000000000000111001",
		b"0000000000000000110111",
		b"0000000000000000110101",
		b"0000000000000000110011",
		b"0000000000000000110001",
		b"0000000000000000101111",
		b"0000000000000000101110",
		b"0000000000000000101100",
		b"0000000000000000101010",
		b"0000000000000000101001",
		b"0000000000000000100111",
		b"0000000000000000100110",
		b"0000000000000000100100",
		b"0000000000000000100011",
		b"0000000000000000100010",
		b"0000000000000000100000",
		b"0000000000000000011111",
		b"0000000000000000011110",
		b"0000000000000000011101",
		b"0000000000000000011100",
		b"0000000000000000011010",
		b"0000000000000000011001",
		b"0000000000000000011000",
		b"0000000000000000010111",
		b"0000000000000000010110",
		b"0000000000000000010101",
		b"0000000000000000010100",
		b"0000000000000000010100",
		b"0000000000000000010011",
		b"0000000000000000010010",
		b"0000000000000000010001",
		b"0000000000000000010000",
		b"0000000000000000010000",
		b"0000000000000000001111",
		b"0000000000000000001110",
		b"0000000000000000001110",
		b"0000000000000000001101",
		b"0000000000000000001100",
		b"0000000000000000001100",
		b"0000000000000000001011",
		b"0000000000000000001011",
		b"0000000000000000001010",
		b"0000000000000000001010",
		b"0000000000000000001001",
		b"0000000000000000001001",
		b"0000000000000000001000",
		b"0000000000000000001000",
		b"0000000000000000000111",
		b"0000000000000000000111",
		b"0000000000000000000111",
		b"0000000000000000000110",
		b"0000000000000000000110",
		b"0000000000000000000101",
		b"0000000000000000000101",
		b"0000000000000000000101",
		b"0000000000000000000101",
		b"0000000000000000000100",
		b"0000000000000000000100",
		b"0000000000000000000100",
		b"0000000000000000000100",
		b"0000000000000000000011",
		b"0000000000000000000011",
		b"0000000000000000000011",
		b"0000000000000000000011",
		b"0000000000000000000011",
		b"0000000000000000000010",
		b"0000000000000000000010",
		b"0000000000000000000010",
		b"0000000000000000000010",
		b"0000000000000000000010",
		b"0000000000000000000010",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000"
	);

end src_rom_pkg;