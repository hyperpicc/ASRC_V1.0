library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package src_rom_pkg is

	constant COE_WIDTH	: integer := 22;
	constant COE_CENTRE	: signed( 21 downto 0 ) := b"0111111101011100001010";

	type COE_ROM_TYPE is array( 4095 downto 0 ) of signed( 21 downto 0 );
	constant COE_ROM	 : COE_ROM_TYPE := (
		b"0111111101011001000111",
		b"0111111101001111111101",
		b"0111111101000000101101",
		b"0111111100101011010111",
		b"0111111100001111111011",
		b"0111111011101110011010",
		b"0111111011000110110101",
		b"0111111010011001001100",
		b"0111111001100101100001",
		b"0111111000101011110101",
		b"0111110111101100001001",
		b"0111110110100110011110",
		b"0111110101011010110110",
		b"0111110100001001010011",
		b"0111110010110001110101",
		b"0111110001010100100000",
		b"0111101111110001010101",
		b"0111101110001000010110",
		b"0111101100011001100110",
		b"0111101010100101000110",
		b"0111101000101010111011",
		b"0111100110101011000101",
		b"0111100100100101101000",
		b"0111100010011010100110",
		b"0111100000001010000100",
		b"0111011101110100000011",
		b"0111011011011000100111",
		b"0111011000110111110011",
		b"0111010110010001101100",
		b"0111010011100110010011",
		b"0111010000110101101110",
		b"0111001110000000000000",
		b"0111001011000101001100",
		b"0111001000000101010111",
		b"0111000101000000100100",
		b"0111000001110110111001",
		b"0110111110101000011001",
		b"0110111011010101001001",
		b"0110110111111101001100",
		b"0110110100100000101001",
		b"0110110000111111100011",
		b"0110101101011010000000",
		b"0110101001110000000011",
		b"0110100110000001110011",
		b"0110100010001111010100",
		b"0110011110011000101011",
		b"0110011010011101111101",
		b"0110010110011111010000",
		b"0110010010011100101010",
		b"0110001110010110001110",
		b"0110001010001100000100",
		b"0110000101111110010001",
		b"0110000001101100111010",
		b"0101111101011000000101",
		b"0101111000111111111000",
		b"0101110100100100011000",
		b"0101110000000101101101",
		b"0101101011100011111010",
		b"0101100110111111001000",
		b"0101100010010111011011",
		b"0101011101101100111001",
		b"0101011000111111101010",
		b"0101010100001111110011",
		b"0101001111011101011010",
		b"0101001010101000100110",
		b"0101000101110001011101",
		b"0101000000111000000110",
		b"0100111011111100100111",
		b"0100110110111111000101",
		b"0100110001111111101001",
		b"0100101100111110011000",
		b"0100100111111011011001",
		b"0100100010110110110010",
		b"0100011101110000101010",
		b"0100011000101001000111",
		b"0100010011100000010001",
		b"0100001110010110001101",
		b"0100001001001011000011",
		b"0100000011111110111000",
		b"0011111110110001110100",
		b"0011111001100011111101",
		b"0011110100010101011010",
		b"0011101111000110010001",
		b"0011101001110110101001",
		b"0011100100100110101000",
		b"0011011111010110010110",
		b"0011011010000101111000",
		b"0011010100110101010101",
		b"0011001111100100110101",
		b"0011001010010100011100",
		b"0011000101000100010010",
		b"0010111111110100011101",
		b"0010111010100101000100",
		b"0010110101010110001101",
		b"0010110000000111111110",
		b"0010101010111010011110",
		b"0010100101101101110011",
		b"0010100000100010000011",
		b"0010011011010111010100",
		b"0010010110001101101101",
		b"0010010001000101010011",
		b"0010001011111110001101",
		b"0010000110111000100001",
		b"0010000001110100010100",
		b"0001111100110001101101",
		b"0001110111110000110001",
		b"0001110010110001100110",
		b"0001101101110100010010",
		b"0001101000111000111010",
		b"0001100011111111100100",
		b"0001011111001000010110",
		b"0001011010010011010100",
		b"0001010101100000100101",
		b"0001010000110000001110",
		b"0001001100000010010011",
		b"0001000111010110111010",
		b"0001000010101110001000",
		b"0000111110001000000001",
		b"0000111001100100101100",
		b"0000110101000100001100",
		b"0000110000100110100110",
		b"0000101100001011111111",
		b"0000100111110100011011",
		b"0000100011011111111111",
		b"0000011111001110101111",
		b"0000011011000000110000",
		b"0000010110110110000101",
		b"0000010010101110110011",
		b"0000001110101010111101",
		b"0000001010101010101000",
		b"0000000110101101110110",
		b"0000000010110100101101",
		b"1111111110111111001111",
		b"1111111011001101011111",
		b"1111110111011111100010",
		b"1111110011110101011010",
		b"1111110000001111001010",
		b"1111101100101100110110",
		b"1111101001001110100000",
		b"1111100101110100001011",
		b"1111100010011101111010",
		b"1111011111001011110000",
		b"1111011011111101101110",
		b"1111011000110011111000",
		b"1111010101101110001111",
		b"1111010010101100110101",
		b"1111001111101111101101",
		b"1111001100110110111001",
		b"1111001010000010011010",
		b"1111000111010010010010",
		b"1111000100100110100010",
		b"1111000001111111001100",
		b"1110111111011100010001",
		b"1110111100111101110011",
		b"1110111010100011110010",
		b"1110111000001110010000",
		b"1110110101111101001101",
		b"1110110011110000101011",
		b"1110110001101000101001",
		b"1110101111100101001000",
		b"1110101101100110001001",
		b"1110101011101011101011",
		b"1110101001110101110000",
		b"1110101000000100010111",
		b"1110100110010111100000",
		b"1110100100101111001011",
		b"1110100011001011011000",
		b"1110100001101100000110",
		b"1110100000010001010100",
		b"1110011110111011000011",
		b"1110011101101001010001",
		b"1110011100011011111110",
		b"1110011011010011001001",
		b"1110011010001110110000",
		b"1110011001001110110010",
		b"1110011000010011001111",
		b"1110010111011100000100",
		b"1110010110101001010001",
		b"1110010101111010110100",
		b"1110010101010000101011",
		b"1110010100101010110100",
		b"1110010100001001001110",
		b"1110010011101011110111",
		b"1110010011010010101100",
		b"1110010010111101101011",
		b"1110010010101100110010",
		b"1110010010100000000000",
		b"1110010010010111010000",
		b"1110010010010010100010",
		b"1110010010010001110001",
		b"1110010010010100111100",
		b"1110010010011100000000",
		b"1110010010100110111010",
		b"1110010010110101100111",
		b"1110010011001000000100",
		b"1110010011011110001101",
		b"1110010011111000000000",
		b"1110010100010101011010",
		b"1110010100110110010111",
		b"1110010101011010110011",
		b"1110010110000010101100",
		b"1110010110101101111110",
		b"1110010111011100100100",
		b"1110011000001110011100",
		b"1110011001000011100010",
		b"1110011001111011110010",
		b"1110011010110111001000",
		b"1110011011110101100000",
		b"1110011100110110110111",
		b"1110011101111011000111",
		b"1110011111000010001110",
		b"1110100000001100000111",
		b"1110100001011000101110",
		b"1110100010100111111111",
		b"1110100011111001110101",
		b"1110100101001110001101",
		b"1110100110100101000001",
		b"1110100111111110001110",
		b"1110101001011001110000",
		b"1110101010110111100001",
		b"1110101100010111011101",
		b"1110101101111001100001",
		b"1110101111011101100110",
		b"1110110001000011101010",
		b"1110110010101011100111",
		b"1110110100010101011000",
		b"1110110110000000111010",
		b"1110110111101110001000",
		b"1110111001011100111100",
		b"1110111011001101010011",
		b"1110111100111111000111",
		b"1110111110110010010101",
		b"1111000000100110110110",
		b"1111000010011100101000",
		b"1111000100010011100101",
		b"1111000110001011101000",
		b"1111001000000100101110",
		b"1111001001111110110000",
		b"1111001011111001101011",
		b"1111001101110101011010",
		b"1111001111110001111001",
		b"1111010001101111000010",
		b"1111010011101100110001",
		b"1111010101101011000010",
		b"1111010111101001110001",
		b"1111011001101000111000",
		b"1111011011101000010011",
		b"1111011101100111111101",
		b"1111011111100111110011",
		b"1111100001100111110000",
		b"1111100011100111101111",
		b"1111100101100111101100",
		b"1111100111100111100011",
		b"1111101001100111001111",
		b"1111101011100110101101",
		b"1111101101100101111000",
		b"1111101111100100101011",
		b"1111110001100011000100",
		b"1111110011100000111101",
		b"1111110101011110010010",
		b"1111110111011011000001",
		b"1111111001010111000100",
		b"1111111011010010011000",
		b"1111111101001100111001",
		b"1111111111000110100100",
		b"0000000000111111010100",
		b"0000000010110111000110",
		b"0000000100101101110110",
		b"0000000110100011100001",
		b"0000001000011000000011",
		b"0000001010001011011010",
		b"0000001011111101100001",
		b"0000001101101110010101",
		b"0000001111011101110011",
		b"0000010001001011111000",
		b"0000010010111000100000",
		b"0000010100100011101010",
		b"0000010110001101010001",
		b"0000010111110101010100",
		b"0000011001011011101110",
		b"0000011011000000011110",
		b"0000011100100011100000",
		b"0000011110000100110010",
		b"0000011111100100010011",
		b"0000100001000001111110",
		b"0000100010011101110010",
		b"0000100011110111101101",
		b"0000100101001111101100",
		b"0000100110100101101101",
		b"0000100111111001101110",
		b"0000101001001011101101",
		b"0000101010011011101001",
		b"0000101011101001011111",
		b"0000101100110101001110",
		b"0000101101111110110100",
		b"0000101111000110010000",
		b"0000110000001011011111",
		b"0000110001001110100001",
		b"0000110010001111010101",
		b"0000110011001101111001",
		b"0000110100001010001011",
		b"0000110101000100001100",
		b"0000110101111011111001",
		b"0000110110110001010010",
		b"0000110111100100010110",
		b"0000111000010101000101",
		b"0000111001000011011101",
		b"0000111001101111011111",
		b"0000111010011001001001",
		b"0000111011000000011011",
		b"0000111011100101010110",
		b"0000111100000111111000",
		b"0000111100101000000001",
		b"0000111101000101110010",
		b"0000111101100001001010",
		b"0000111101111010001010",
		b"0000111110010000110001",
		b"0000111110100101000000",
		b"0000111110110110110111",
		b"0000111111000110010110",
		b"0000111111010011011111",
		b"0000111111011110010000",
		b"0000111111100110101100",
		b"0000111111101100110011",
		b"0000111111110000100101",
		b"0000111111110010000100",
		b"0000111111110001010000",
		b"0000111111101110001010",
		b"0000111111101000110011",
		b"0000111111100001001100",
		b"0000111111010111010111",
		b"0000111111001011010101",
		b"0000111110111101000111",
		b"0000111110101100101110",
		b"0000111110011010001101",
		b"0000111110000101100011",
		b"0000111101101110110100",
		b"0000111101010110000000",
		b"0000111100111011001010",
		b"0000111100011110010010",
		b"0000111011111111011100",
		b"0000111011011110101000",
		b"0000111010111011111001",
		b"0000111010010111010000",
		b"0000111001110000110000",
		b"0000111001001000011010",
		b"0000111000011110010010",
		b"0000110111110010011000",
		b"0000110111000100101111",
		b"0000110110010101011010",
		b"0000110101100100011011",
		b"0000110100110001110100",
		b"0000110011111101100111",
		b"0000110011000111110111",
		b"0000110010010000100110",
		b"0000110001010111110111",
		b"0000110000011101101101",
		b"0000101111100010001010",
		b"0000101110100101010000",
		b"0000101101100111000010",
		b"0000101100100111100011",
		b"0000101011100110110110",
		b"0000101010100100111101",
		b"0000101001100001111100",
		b"0000101000011101110100",
		b"0000100111011000101000",
		b"0000100110010010011100",
		b"0000100101001011010010",
		b"0000100100000011001101",
		b"0000100010111010010000",
		b"0000100001110000011110",
		b"0000100000100101111010",
		b"0000011111011010100110",
		b"0000011110001110100110",
		b"0000011101000001111100",
		b"0000011011110100101011",
		b"0000011010100110110110",
		b"0000011001011000100001",
		b"0000011000001001101110",
		b"0000010110111010011111",
		b"0000010101101010111001",
		b"0000010100011010111101",
		b"0000010011001010101111",
		b"0000010001111010010010",
		b"0000010000101001101001",
		b"0000001111011000110110",
		b"0000001110000111111100",
		b"0000001100110110111110",
		b"0000001011100110000000",
		b"0000001010010101000011",
		b"0000001001000100001011",
		b"0000000111110011011011",
		b"0000000110100010110101",
		b"0000000101010010011100",
		b"0000000100000010010011",
		b"0000000010110010011101",
		b"0000000001100010111100",
		b"0000000000010011110011",
		b"1111111111000101000100",
		b"1111111101110110110011",
		b"1111111100101001000001",
		b"1111111011011011110010",
		b"1111111010001111001000",
		b"1111111001000011000101",
		b"1111110111110111101100",
		b"1111110110101100111111",
		b"1111110101100011000001",
		b"1111110100011001110011",
		b"1111110011010001011001",
		b"1111110010001001110101",
		b"1111110001000011001001",
		b"1111101111111101010110",
		b"1111101110111000100000",
		b"1111101101110100101000",
		b"1111101100110001110000",
		b"1111101011101111111011",
		b"1111101010101111001010",
		b"1111101001101111011111",
		b"1111101000110000111100",
		b"1111100111110011100011",
		b"1111100110110111010110",
		b"1111100101111100010110",
		b"1111100101000010100110",
		b"1111100100001010000110",
		b"1111100011010010111000",
		b"1111100010011100111110",
		b"1111100001101000011010",
		b"1111100000110101001100",
		b"1111100000000011010111",
		b"1111011111010010111010",
		b"1111011110100011111001",
		b"1111011101110110010011",
		b"1111011101001010001010",
		b"1111011100011111011111",
		b"1111011011110110010100",
		b"1111011011001110101000",
		b"1111011010101000011101",
		b"1111011010000011110101",
		b"1111011001100000101110",
		b"1111011000111111001100",
		b"1111011000011111001101",
		b"1111011000000000110011",
		b"1111010111100011111110",
		b"1111010111001000110000",
		b"1111010110101111000111",
		b"1111010110010111000101",
		b"1111010110000000101010",
		b"1111010101101011110110",
		b"1111010101011000101010",
		b"1111010101000111000110",
		b"1111010100110111001001",
		b"1111010100101000110100",
		b"1111010100011100001000",
		b"1111010100010001000010",
		b"1111010100000111100101",
		b"1111010011111111101111",
		b"1111010011111001100001",
		b"1111010011110100111001",
		b"1111010011110001111000",
		b"1111010011110000011110",
		b"1111010011110000101001",
		b"1111010011110010011010",
		b"1111010011110101101111",
		b"1111010011111010101001",
		b"1111010100000001000110",
		b"1111010100001001000111",
		b"1111010100010010101001",
		b"1111010100011101101101",
		b"1111010100101010010001",
		b"1111010100111000010101",
		b"1111010101000111110111",
		b"1111010101011000110111",
		b"1111010101101011010100",
		b"1111010101111111001100",
		b"1111010110010100011111",
		b"1111010110101011001011",
		b"1111010111000011001111",
		b"1111010111011100101001",
		b"1111010111110111011001",
		b"1111011000010011011110",
		b"1111011000110000110101",
		b"1111011001001111011101",
		b"1111011001101111010101",
		b"1111011010010000011011",
		b"1111011010110010101111",
		b"1111011011010110001101",
		b"1111011011111010110101",
		b"1111011100100000100110",
		b"1111011101000111011100",
		b"1111011101101111011000",
		b"1111011110011000010110",
		b"1111011111000010010101",
		b"1111011111101101010100",
		b"1111100000011001010001",
		b"1111100001000110001001",
		b"1111100001110011111011",
		b"1111100010100010100101",
		b"1111100011010010000110",
		b"1111100100000010011010",
		b"1111100100110011100001",
		b"1111100101100101011000",
		b"1111100110010111111110",
		b"1111100111001011010000",
		b"1111100111111111001100",
		b"1111101000110011110000",
		b"1111101001101000111011",
		b"1111101010011110101010",
		b"1111101011010100111011",
		b"1111101100001011101100",
		b"1111101101000010111011",
		b"1111101101111010100110",
		b"1111101110110010101011",
		b"1111101111101011001000",
		b"1111110000100011111010",
		b"1111110001011101000000",
		b"1111110010010110010111",
		b"1111110011001111111110",
		b"1111110100001001110001",
		b"1111110101000011110000",
		b"1111110101111101111000",
		b"1111110110111000000110",
		b"1111110111110010011001",
		b"1111111000101100110000",
		b"1111111001100111000110",
		b"1111111010100001011011",
		b"1111111011011011101101",
		b"1111111100010101111001",
		b"1111111101001111111110",
		b"1111111110001001111001",
		b"1111111111000011101001",
		b"1111111111111101001010",
		b"0000000000110110011100",
		b"0000000001101111011101",
		b"0000000010101000001010",
		b"0000000011100000100010",
		b"0000000100011000100010",
		b"0000000101010000001001",
		b"0000000110000111010101",
		b"0000000110111110000100",
		b"0000000111110100010101",
		b"0000001000101010000101",
		b"0000001001011111010010",
		b"0000001010010011111011",
		b"0000001011000111111111",
		b"0000001011111011011011",
		b"0000001100101110001110",
		b"0000001101100000010111",
		b"0000001110010001110011",
		b"0000001111000010100001",
		b"0000001111110010011111",
		b"0000010000100001101101",
		b"0000010001010000001000",
		b"0000010001111101110000",
		b"0000010010101010100010",
		b"0000010011010110011101",
		b"0000010100000001100001",
		b"0000010100101011101011",
		b"0000010101010100111011",
		b"0000010101111101001111",
		b"0000010110100100100110",
		b"0000010111001010111111",
		b"0000010111110000011001",
		b"0000011000010100110011",
		b"0000011000111000001011",
		b"0000011001011010100001",
		b"0000011001111011110100",
		b"0000011010011100000010",
		b"0000011010111011001100",
		b"0000011011011001010000",
		b"0000011011110110001101",
		b"0000011100010010000011",
		b"0000011100101100110001",
		b"0000011101000110010110",
		b"0000011101011110110010",
		b"0000011101110110000100",
		b"0000011110001100001100",
		b"0000011110100001001001",
		b"0000011110110100111010",
		b"0000011111000111100000",
		b"0000011111011000111001",
		b"0000011111101001000110",
		b"0000011111111000000111",
		b"0000100000000101111010",
		b"0000100000010010100001",
		b"0000100000011101111010",
		b"0000100000101000000110",
		b"0000100000110001000101",
		b"0000100000111000110110",
		b"0000100000111111011001",
		b"0000100001000100110000",
		b"0000100001001000111001",
		b"0000100001001011110101",
		b"0000100001001101100101",
		b"0000100001001110001000",
		b"0000100001001101011110",
		b"0000100001001011101001",
		b"0000100001001000101000",
		b"0000100001000100011100",
		b"0000100000111111000101",
		b"0000100000111000100011",
		b"0000100000110000111000",
		b"0000100000101000000100",
		b"0000100000011110000111",
		b"0000100000010011000011",
		b"0000100000000110110111",
		b"0000011111111001100100",
		b"0000011111101011001011",
		b"0000011111011011101110",
		b"0000011111001011001100",
		b"0000011110111001100111",
		b"0000011110100110111111",
		b"0000011110010011010110",
		b"0000011101111110101100",
		b"0000011101101001000011",
		b"0000011101010010011011",
		b"0000011100111010110101",
		b"0000011100100010010011",
		b"0000011100001000110101",
		b"0000011011101110011101",
		b"0000011011010011001100",
		b"0000011010110111000011",
		b"0000011010011010000011",
		b"0000011001111100001110",
		b"0000011001011101100101",
		b"0000011000111110001000",
		b"0000011000011101111011",
		b"0000010111111100111100",
		b"0000010111011011001111",
		b"0000010110111000110100",
		b"0000010110010101101110",
		b"0000010101110001111100",
		b"0000010101001101100001",
		b"0000010100101000011110",
		b"0000010100000010110101",
		b"0000010011011100100111",
		b"0000010010110101110110",
		b"0000010010001110100011",
		b"0000010001100110101111",
		b"0000010000111110011100",
		b"0000010000010101101101",
		b"0000001111101100100001",
		b"0000001111000010111011",
		b"0000001110011000111101",
		b"0000001101101110101000",
		b"0000001101000011111101",
		b"0000001100011000111111",
		b"0000001011101101101110",
		b"0000001011000010001101",
		b"0000001010010110011100",
		b"0000001001101010011111",
		b"0000001000111110010101",
		b"0000001000010010000010",
		b"0000000111100101100110",
		b"0000000110111001000011",
		b"0000000110001100011010",
		b"0000000101011111101110",
		b"0000000100110011000000",
		b"0000000100000110010010",
		b"0000000011011001100100",
		b"0000000010101100111001",
		b"0000000010000000010011",
		b"0000000001010011110010",
		b"0000000000100111011000",
		b"1111111111111011001000",
		b"1111111111001111000010",
		b"1111111110100011001000",
		b"1111111101110111011100",
		b"1111111101001011111110",
		b"1111111100100000110001",
		b"1111111011110101110111",
		b"1111111011001011001111",
		b"1111111010100000111101",
		b"1111111001110111000001",
		b"1111111001001101011100",
		b"1111111000100100010001",
		b"1111110111111011100001",
		b"1111110111010011001100",
		b"1111110110101011010100",
		b"1111110110000011111011",
		b"1111110101011101000010",
		b"1111110100110110101010",
		b"1111110100010000110100",
		b"1111110011101011100010",
		b"1111110011000110110101",
		b"1111110010100010101101",
		b"1111110001111111001101",
		b"1111110001011100010101",
		b"1111110000111010000110",
		b"1111110000011000100001",
		b"1111101111110111101000",
		b"1111101111010111011100",
		b"1111101110110111111101",
		b"1111101110011001001100",
		b"1111101101111011001010",
		b"1111101101011101111001",
		b"1111101101000001011001",
		b"1111101100100101101011",
		b"1111101100001010110000",
		b"1111101011110000101000",
		b"1111101011010111010100",
		b"1111101010111110110101",
		b"1111101010100111001100",
		b"1111101010010000011010",
		b"1111101001111010011110",
		b"1111101001100101011010",
		b"1111101001010001001110",
		b"1111101000111101111011",
		b"1111101000101011100000",
		b"1111101000011010000000",
		b"1111101000001001011001",
		b"1111100111111001101100",
		b"1111100111101010111011",
		b"1111100111011101000100",
		b"1111100111010000001001",
		b"1111100111000100001001",
		b"1111100110111001000101",
		b"1111100110101110111101",
		b"1111100110100101110010",
		b"1111100110011101100010",
		b"1111100110010110001111",
		b"1111100110001111111000",
		b"1111100110001010011110",
		b"1111100110000110000000",
		b"1111100110000010011110",
		b"1111100101111111111001",
		b"1111100101111110010000",
		b"1111100101111101100011",
		b"1111100101111101110001",
		b"1111100101111110111100",
		b"1111100110000001000001",
		b"1111100110000100000010",
		b"1111100110000111111110",
		b"1111100110001100110011",
		b"1111100110010010100011",
		b"1111100110011001001101",
		b"1111100110100000110000",
		b"1111100110101001001011",
		b"1111100110110010011111",
		b"1111100110111100101011",
		b"1111100111000111101101",
		b"1111100111010011100111",
		b"1111100111100000010110",
		b"1111100111101101111011",
		b"1111100111111100010100",
		b"1111101000001011100010",
		b"1111101000011011100010",
		b"1111101000101100010101",
		b"1111101000111101111010",
		b"1111101001010000010000",
		b"1111101001100011010110",
		b"1111101001110111001011",
		b"1111101010001011101111",
		b"1111101010100001000000",
		b"1111101010110110111110",
		b"1111101011001101101000",
		b"1111101011100100111100",
		b"1111101011111100111010",
		b"1111101100010101100001",
		b"1111101100101110110000",
		b"1111101101001000100101",
		b"1111101101100011000001",
		b"1111101101111110000000",
		b"1111101110011001100011",
		b"1111101110110101101001",
		b"1111101111010010010000",
		b"1111101111101111010111",
		b"1111110000001100111101",
		b"1111110000101011000001",
		b"1111110001001001100010",
		b"1111110001101000011110",
		b"1111110010000111110101",
		b"1111110010100111100100",
		b"1111110011000111101100",
		b"1111110011101000001010",
		b"1111110100001000111110",
		b"1111110100101010000101",
		b"1111110101001011100000",
		b"1111110101101101001101",
		b"1111110110001111001010",
		b"1111110110110001010110",
		b"1111110111010011110000",
		b"1111110111110110010110",
		b"1111111000011001001000",
		b"1111111000111100000101",
		b"1111111001011111001001",
		b"1111111010000010010110",
		b"1111111010100101101000",
		b"1111111011001001000000",
		b"1111111011101100011011",
		b"1111111100001111111001",
		b"1111111100110011011000",
		b"1111111101010110110111",
		b"1111111101111010010100",
		b"1111111110011101101111",
		b"1111111111000001000110",
		b"1111111111100100010111",
		b"0000000000000111100010",
		b"0000000000101010100110",
		b"0000000001001101100001",
		b"0000000001110000010001",
		b"0000000010010010110111",
		b"0000000010110101010000",
		b"0000000011010111011011",
		b"0000000011111001010111",
		b"0000000100011011000100",
		b"0000000100111100011111",
		b"0000000101011101101000",
		b"0000000101111110011110",
		b"0000000110011110111111",
		b"0000000110111111001010",
		b"0000000111011110111111",
		b"0000000111111110011100",
		b"0000001000011101100001",
		b"0000001000111100001011",
		b"0000001001011010011011",
		b"0000001001111000001111",
		b"0000001010010101100110",
		b"0000001010110010011111",
		b"0000001011001110111010",
		b"0000001011101010110101",
		b"0000001100000110001111",
		b"0000001100100001001000",
		b"0000001100111011100000",
		b"0000001101010101010011",
		b"0000001101101110100100",
		b"0000001110000111001111",
		b"0000001110011111010101",
		b"0000001110110110110101",
		b"0000001111001101101110",
		b"0000001111100100000000",
		b"0000001111111001101001",
		b"0000010000001110101010",
		b"0000010000100011000001",
		b"0000010000110110101110",
		b"0000010001001001110001",
		b"0000010001011100001000",
		b"0000010001101101110011",
		b"0000010001111110110011",
		b"0000010010001111000110",
		b"0000010010011110101011",
		b"0000010010101101100011",
		b"0000010010111011101110",
		b"0000010011001001001010",
		b"0000010011010101110111",
		b"0000010011100001110110",
		b"0000010011101101000101",
		b"0000010011110111100101",
		b"0000010100000001010110",
		b"0000010100001010010110",
		b"0000010100010010100111",
		b"0000010100011010001000",
		b"0000010100100000111000",
		b"0000010100100110111000",
		b"0000010100101100000111",
		b"0000010100110000100110",
		b"0000010100110100010101",
		b"0000010100110111010011",
		b"0000010100111001100001",
		b"0000010100111010111110",
		b"0000010100111011101100",
		b"0000010100111011101001",
		b"0000010100111010110110",
		b"0000010100111001010100",
		b"0000010100110111000010",
		b"0000010100110100000001",
		b"0000010100110000010001",
		b"0000010100101011110010",
		b"0000010100100110100100",
		b"0000010100100000101001",
		b"0000010100011001111111",
		b"0000010100010010101001",
		b"0000010100001010100101",
		b"0000010100000001110101",
		b"0000010011111000011000",
		b"0000010011101110010000",
		b"0000010011100011011101",
		b"0000010011010111111111",
		b"0000010011001011110111",
		b"0000010010111111000110",
		b"0000010010110001101100",
		b"0000010010100011101001",
		b"0000010010010100111111",
		b"0000010010000101101110",
		b"0000010001110101110110",
		b"0000010001100101011001",
		b"0000010001010100010110",
		b"0000010001000010110000",
		b"0000010000110000100110",
		b"0000010000011101111001",
		b"0000010000001010101010",
		b"0000001111110110111010",
		b"0000001111100010101010",
		b"0000001111001101111010",
		b"0000001110111000101011",
		b"0000001110100010111110",
		b"0000001110001100110101",
		b"0000001101110110001111",
		b"0000001101011111001110",
		b"0000001101000111110011",
		b"0000001100101111111110",
		b"0000001100010111110001",
		b"0000001011111111001101",
		b"0000001011100110010001",
		b"0000001011001101000000",
		b"0000001010110011011011",
		b"0000001010011001100001",
		b"0000001001111111010110",
		b"0000001001100100111000",
		b"0000001001001010001001",
		b"0000001000101111001011",
		b"0000001000010011111111",
		b"0000000111111000100100",
		b"0000000111011100111101",
		b"0000000111000001001010",
		b"0000000110100101001101",
		b"0000000110001001000110",
		b"0000000101101100110110",
		b"0000000101010000011111",
		b"0000000100110100000010",
		b"0000000100010111011111",
		b"0000000011111010110111",
		b"0000000011011110001100",
		b"0000000011000001011111",
		b"0000000010100100110001",
		b"0000000010001000000010",
		b"0000000001101011010100",
		b"0000000001001110101000",
		b"0000000000110001111111",
		b"0000000000010101011001",
		b"1111111111111000111000",
		b"1111111111011100011101",
		b"1111111111000000001001",
		b"1111111110100011111101",
		b"1111111110000111111001",
		b"1111111101101011111111",
		b"1111111101010000010000",
		b"1111111100110100101100",
		b"1111111100011001010110",
		b"1111111011111110001100",
		b"1111111011100011010001",
		b"1111111011001000100110",
		b"1111111010101110001011",
		b"1111111010010100000001",
		b"1111111001111010001001",
		b"1111111001100000100100",
		b"1111111001000111010011",
		b"1111111000101110010111",
		b"1111111000010101110000",
		b"1111110111111101011111",
		b"1111110111100101100101",
		b"1111110111001110000100",
		b"1111110110110110111010",
		b"1111110110100000001011",
		b"1111110110001001110101",
		b"1111110101110011111010",
		b"1111110101011110011011",
		b"1111110101001001011000",
		b"1111110100110100110010",
		b"1111110100100000101001",
		b"1111110100001100111111",
		b"1111110011111001110011",
		b"1111110011100111000111",
		b"1111110011010100111010",
		b"1111110011000011001111",
		b"1111110010110010000100",
		b"1111110010100001011010",
		b"1111110010010001010011",
		b"1111110010000001101110",
		b"1111110001110010101100",
		b"1111110001100100001110",
		b"1111110001010110010011",
		b"1111110001001000111101",
		b"1111110000111100001011",
		b"1111110000101111111110",
		b"1111110000100100010110",
		b"1111110000011001010100",
		b"1111110000001110110111",
		b"1111110000000101000001",
		b"1111101111111011110001",
		b"1111101111110011000111",
		b"1111101111101011000101",
		b"1111101111100011101001",
		b"1111101111011100110100",
		b"1111101111010110100110",
		b"1111101111010000111111",
		b"1111101111001100000000",
		b"1111101111000111101000",
		b"1111101111000011111000",
		b"1111101111000000101111",
		b"1111101110111110001110",
		b"1111101110111100010100",
		b"1111101110111011000001",
		b"1111101110111010010110",
		b"1111101110111010010010",
		b"1111101110111010110101",
		b"1111101110111011111111",
		b"1111101110111101110000",
		b"1111101111000000000111",
		b"1111101111000011000101",
		b"1111101111000110101001",
		b"1111101111001010110011",
		b"1111101111001111100011",
		b"1111101111010100111000",
		b"1111101111011010110011",
		b"1111101111100001010010",
		b"1111101111101000010101",
		b"1111101111101111111101",
		b"1111101111111000001000",
		b"1111110000000000110111",
		b"1111110000001010001001",
		b"1111110000010011111101",
		b"1111110000011110010011",
		b"1111110000101001001011",
		b"1111110000110100100011",
		b"1111110001000000011101",
		b"1111110001001100110110",
		b"1111110001011001101111",
		b"1111110001100111000111",
		b"1111110001110100111101",
		b"1111110010000011010001",
		b"1111110010010010000010",
		b"1111110010100001010000",
		b"1111110010110000111010",
		b"1111110011000000111111",
		b"1111110011010001011111",
		b"1111110011100010011000",
		b"1111110011110011101100",
		b"1111110100000101010111",
		b"1111110100010111011011",
		b"1111110100101001110110",
		b"1111110100111100100111",
		b"1111110101001111101110",
		b"1111110101100011001010",
		b"1111110101110110111011",
		b"1111110110001010111110",
		b"1111110110011111010101",
		b"1111110110110011111101",
		b"1111110111001000110111",
		b"1111110111011110000001",
		b"1111110111110011011010",
		b"1111111000001001000011",
		b"1111111000011110111001",
		b"1111111000110100111100",
		b"1111111001001011001011",
		b"1111111001100001100110",
		b"1111111001111000001100",
		b"1111111010001110111011",
		b"1111111010100101110100",
		b"1111111010111100110100",
		b"1111111011010011111100",
		b"1111111011101011001010",
		b"1111111100000010011101",
		b"1111111100011001110101",
		b"1111111100110001010010",
		b"1111111101001000110001",
		b"1111111101100000010010",
		b"1111111101110111110101",
		b"1111111110001111011000",
		b"1111111110100110111010",
		b"1111111110111110011100",
		b"1111111111010101111100",
		b"1111111111101101011000",
		b"0000000000000100110001",
		b"0000000000011100000101",
		b"0000000000110011010101",
		b"0000000001001010011101",
		b"0000000001100001011111",
		b"0000000001111000011010",
		b"0000000010001111001011",
		b"0000000010100101110011",
		b"0000000010111100010010",
		b"0000000011010010100101",
		b"0000000011101000101101",
		b"0000000011111110101000",
		b"0000000100010100010110",
		b"0000000100101001110110",
		b"0000000100111111000111",
		b"0000000101010100001001",
		b"0000000101101000111100",
		b"0000000101111101011101",
		b"0000000110010001101101",
		b"0000000110100101101011",
		b"0000000110111001010110",
		b"0000000111001100101110",
		b"0000000111011111110001",
		b"0000000111110010100000",
		b"0000001000000100111010",
		b"0000001000010110111110",
		b"0000001000101000101011",
		b"0000001000111010000010",
		b"0000001001001011000000",
		b"0000001001011011100111",
		b"0000001001101011110101",
		b"0000001001111011101010",
		b"0000001010001011000110",
		b"0000001010011010000111",
		b"0000001010101000101110",
		b"0000001010110110111001",
		b"0000001011000100101010",
		b"0000001011010001111110",
		b"0000001011011110110110",
		b"0000001011101011010010",
		b"0000001011110111010001",
		b"0000001100000010110010",
		b"0000001100001101110110",
		b"0000001100011000011011",
		b"0000001100100010100011",
		b"0000001100101100001100",
		b"0000001100110101010110",
		b"0000001100111110000001",
		b"0000001101000110001101",
		b"0000001101001101111010",
		b"0000001101010101000111",
		b"0000001101011011110100",
		b"0000001101100010000001",
		b"0000001101100111101110",
		b"0000001101101100111011",
		b"0000001101110001101000",
		b"0000001101110101110100",
		b"0000001101111001100000",
		b"0000001101111100101100",
		b"0000001101111111010111",
		b"0000001110000001100010",
		b"0000001110000011001100",
		b"0000001110000100010110",
		b"0000001110000100111111",
		b"0000001110000101001000",
		b"0000001110000100110001",
		b"0000001110000011111010",
		b"0000001110000010100011",
		b"0000001110000000101100",
		b"0000001101111110010110",
		b"0000001101111011100000",
		b"0000001101111000001010",
		b"0000001101110100010110",
		b"0000001101110000000011",
		b"0000001101101011010001",
		b"0000001101100110000001",
		b"0000001101100000010010",
		b"0000001101011010000110",
		b"0000001101010011011100",
		b"0000001101001100010110",
		b"0000001101000100110010",
		b"0000001100111100110010",
		b"0000001100110100010110",
		b"0000001100101011011110",
		b"0000001100100010001010",
		b"0000001100011000011100",
		b"0000001100001110010011",
		b"0000001100000011110000",
		b"0000001011111000110100",
		b"0000001011101101011110",
		b"0000001011100001110000",
		b"0000001011010101101010",
		b"0000001011001001001100",
		b"0000001010111100010110",
		b"0000001010101111001010",
		b"0000001010100001101000",
		b"0000001010010011110001",
		b"0000001010000101100100",
		b"0000001001110111000011",
		b"0000001001101000001110",
		b"0000001001011001000110",
		b"0000001001001001101011",
		b"0000001000111001111110",
		b"0000001000101001111111",
		b"0000001000011001110000",
		b"0000001000001001010000",
		b"0000000111111000100001",
		b"0000000111100111100011",
		b"0000000111010110010111",
		b"0000000111000100111101",
		b"0000000110110011010101",
		b"0000000110100001100010",
		b"0000000110001111100011",
		b"0000000101111101011001",
		b"0000000101101011000101",
		b"0000000101011000100111",
		b"0000000101000110000000",
		b"0000000100110011010001",
		b"0000000100100000011010",
		b"0000000100001101011100",
		b"0000000011111010011001",
		b"0000000011100111001111",
		b"0000000011010100000001",
		b"0000000011000000101111",
		b"0000000010101101011010",
		b"0000000010011010000010",
		b"0000000010000110101000",
		b"0000000001110011001100",
		b"0000000001011111110001",
		b"0000000001001100010101",
		b"0000000000111000111010",
		b"0000000000100101100000",
		b"0000000000010010001001",
		b"1111111111111110110100",
		b"1111111111101011100100",
		b"1111111111011000010111",
		b"1111111111000101001111",
		b"1111111110110010001101",
		b"1111111110011111010001",
		b"1111111110001100011100",
		b"1111111101111001101110",
		b"1111111101100111001001",
		b"1111111101010100101100",
		b"1111111101000010011001",
		b"1111111100110000010000",
		b"1111111100011110010001",
		b"1111111100001100011110",
		b"1111111011111010110111",
		b"1111111011101001011101",
		b"1111111011011000001111",
		b"1111111011000111001111",
		b"1111111010110110011101",
		b"1111111010100101111011",
		b"1111111010010101100111",
		b"1111111010000101100011",
		b"1111111001110101110000",
		b"1111111001100110001110",
		b"1111111001010110111101",
		b"1111111001000111111110",
		b"1111111000111001010001",
		b"1111111000101010110111",
		b"1111111000011100110001",
		b"1111111000001110111110",
		b"1111111000000001100000",
		b"1111110111110100010110",
		b"1111110111100111100001",
		b"1111110111011011000010",
		b"1111110111001110111001",
		b"1111110111000011000101",
		b"1111110110110111101001",
		b"1111110110101100100011",
		b"1111110110100001110100",
		b"1111110110010111011101",
		b"1111110110001101011110",
		b"1111110110000011110111",
		b"1111110101111010101001",
		b"1111110101110001110011",
		b"1111110101101001010110",
		b"1111110101100001010010",
		b"1111110101011001100111",
		b"1111110101010010010110",
		b"1111110101001011011111",
		b"1111110101000101000010",
		b"1111110100111110111111",
		b"1111110100111001010110",
		b"1111110100110100000111",
		b"1111110100101111010011",
		b"1111110100101010111010",
		b"1111110100100110111011",
		b"1111110100100011010110",
		b"1111110100100000001101",
		b"1111110100011101011110",
		b"1111110100011011001010",
		b"1111110100011001010001",
		b"1111110100010111110011",
		b"1111110100010110110000",
		b"1111110100010110000111",
		b"1111110100010101111001",
		b"1111110100010110000110",
		b"1111110100010110101101",
		b"1111110100010111101111",
		b"1111110100011001001010",
		b"1111110100011011000001",
		b"1111110100011101010001",
		b"1111110100011111111011",
		b"1111110100100010111111",
		b"1111110100100110011101",
		b"1111110100101010010100",
		b"1111110100101110100100",
		b"1111110100110011001101",
		b"1111110100111000001110",
		b"1111110100111101101001",
		b"1111110101000011011011",
		b"1111110101001001100101",
		b"1111110101010000000111",
		b"1111110101010111000000",
		b"1111110101011110010001",
		b"1111110101100101111000",
		b"1111110101101101110101",
		b"1111110101110110001000",
		b"1111110101111110110001",
		b"1111110110000111110000",
		b"1111110110010001000011",
		b"1111110110011010101011",
		b"1111110110100100100111",
		b"1111110110101110110110",
		b"1111110110111001011001",
		b"1111110111000100001111",
		b"1111110111001111010111",
		b"1111110111011010110001",
		b"1111110111100110011101",
		b"1111110111110010011010",
		b"1111110111111110100111",
		b"1111111000001011000100",
		b"1111111000010111110001",
		b"1111111000100100101101",
		b"1111111000110001111000",
		b"1111111000111111010001",
		b"1111111001001100110111",
		b"1111111001011010101011",
		b"1111111001101000101011",
		b"1111111001110110110111",
		b"1111111010000101001110",
		b"1111111010010011110000",
		b"1111111010100010011101",
		b"1111111010110001010100",
		b"1111111011000000010011",
		b"1111111011001111011100",
		b"1111111011011110101100",
		b"1111111011101110000100",
		b"1111111011111101100100",
		b"1111111100001101001001",
		b"1111111100011100110100",
		b"1111111100101100100101",
		b"1111111100111100011010",
		b"1111111101001100010100",
		b"1111111101011100010001",
		b"1111111101101100010001",
		b"1111111101111100010011",
		b"1111111110001100011000",
		b"1111111110011100011101",
		b"1111111110101100100011",
		b"1111111110111100101001",
		b"1111111111001100101111",
		b"1111111111011100110100",
		b"1111111111101100110111",
		b"1111111111111100110111",
		b"0000000000001100110101",
		b"0000000000011100110000",
		b"0000000000101100100111",
		b"0000000000111100011001",
		b"0000000001001100000111",
		b"0000000001011011101110",
		b"0000000001101011010000",
		b"0000000001111010101011",
		b"0000000010001001111111",
		b"0000000010011001001100",
		b"0000000010101000010000",
		b"0000000010110111001011",
		b"0000000011000101111110",
		b"0000000011010100100110",
		b"0000000011100011000101",
		b"0000000011110001011000",
		b"0000000011111111100001",
		b"0000000100001101011110",
		b"0000000100011011001111",
		b"0000000100101000110011",
		b"0000000100110110001010",
		b"0000000101000011010100",
		b"0000000101010000010000",
		b"0000000101011100111110",
		b"0000000101101001011101",
		b"0000000101110101101100",
		b"0000000110000001101101",
		b"0000000110001101011101",
		b"0000000110011000111101",
		b"0000000110100100001101",
		b"0000000110101111001100",
		b"0000000110111001111001",
		b"0000000111000100010101",
		b"0000000111001110011110",
		b"0000000111011000010110",
		b"0000000111100001111010",
		b"0000000111101011001100",
		b"0000000111110100001011",
		b"0000000111111100110110",
		b"0000001000000101001110",
		b"0000001000001101010010",
		b"0000001000010101000010",
		b"0000001000011100011101",
		b"0000001000100011100100",
		b"0000001000101010010110",
		b"0000001000110000110011",
		b"0000001000110110111010",
		b"0000001000111100101101",
		b"0000001001000010001010",
		b"0000001001000111010010",
		b"0000001001001100000100",
		b"0000001001010000100000",
		b"0000001001010100100110",
		b"0000001001011000010111",
		b"0000001001011011110001",
		b"0000001001011110110101",
		b"0000001001100001100011",
		b"0000001001100011111011",
		b"0000001001100101111101",
		b"0000001001100111101000",
		b"0000001001101000111110",
		b"0000001001101001111101",
		b"0000001001101010100110",
		b"0000001001101010111000",
		b"0000001001101010110101",
		b"0000001001101010011100",
		b"0000001001101001101101",
		b"0000001001101000100111",
		b"0000001001100111001101",
		b"0000001001100101011100",
		b"0000001001100011010110",
		b"0000001001100000111011",
		b"0000001001011110001010",
		b"0000001001011011000101",
		b"0000001001010111101010",
		b"0000001001010011111011",
		b"0000001001001111110111",
		b"0000001001001011011111",
		b"0000001001000110110011",
		b"0000001001000001110011",
		b"0000001000111100011111",
		b"0000001000110110111000",
		b"0000001000110000111110",
		b"0000001000101010110000",
		b"0000001000100100010001",
		b"0000001000011101011110",
		b"0000001000010110011010",
		b"0000001000001111000100",
		b"0000001000000111011101",
		b"0000000111111111100100",
		b"0000000111110111011011",
		b"0000000111101111000001",
		b"0000000111100110011000",
		b"0000000111011101011110",
		b"0000000111010100010101",
		b"0000000111001010111101",
		b"0000000111000001010111",
		b"0000000110110111100010",
		b"0000000110101101011111",
		b"0000000110100011001111",
		b"0000000110011000110010",
		b"0000000110001110001000",
		b"0000000110000011010010",
		b"0000000101111000010000",
		b"0000000101101101000010",
		b"0000000101100001101010",
		b"0000000101010110000111",
		b"0000000101001010011010",
		b"0000000100111110100011",
		b"0000000100110010100100",
		b"0000000100100110011011",
		b"0000000100011010001010",
		b"0000000100001101110010",
		b"0000000100000001010010",
		b"0000000011110100101011",
		b"0000000011100111111101",
		b"0000000011011011001010",
		b"0000000011001110010001",
		b"0000000011000001010011",
		b"0000000010110100010001",
		b"0000000010100111001010",
		b"0000000010011010000000",
		b"0000000010001100110011",
		b"0000000001111111100100",
		b"0000000001110010010010",
		b"0000000001100100111110",
		b"0000000001010111101001",
		b"0000000001001010010100",
		b"0000000000111100111110",
		b"0000000000101111101000",
		b"0000000000100010010011",
		b"0000000000010101000000",
		b"0000000000000111101110",
		b"1111111111111010011110",
		b"1111111111101101010001",
		b"1111111111100000000110",
		b"1111111111010011000000",
		b"1111111111000101111101",
		b"1111111110111000111110",
		b"1111111110101100000101",
		b"1111111110011111010000",
		b"1111111110010010100010",
		b"1111111110000101111010",
		b"1111111101111001011000",
		b"1111111101101100111101",
		b"1111111101100000101010",
		b"1111111101010100011111",
		b"1111111101001000011100",
		b"1111111100111100100001",
		b"1111111100110000110000",
		b"1111111100100101001000",
		b"1111111100011001101010",
		b"1111111100001110010110",
		b"1111111100000011001101",
		b"1111111011111000001111",
		b"1111111011101101011101",
		b"1111111011100010110110",
		b"1111111011011000011011",
		b"1111111011001110001100",
		b"1111111011000100001010",
		b"1111111010111010010101",
		b"1111111010110000101110",
		b"1111111010100111010100",
		b"1111111010011110001000",
		b"1111111010010101001010",
		b"1111111010001100011011",
		b"1111111010000011111010",
		b"1111111001111011101001",
		b"1111111001110011100111",
		b"1111111001101011110100",
		b"1111111001100100010001",
		b"1111111001011100111110",
		b"1111111001010101111100",
		b"1111111001001111001001",
		b"1111111001001000101000",
		b"1111111001000010010111",
		b"1111111000111100010111",
		b"1111111000110110101000",
		b"1111111000110001001010",
		b"1111111000101011111110",
		b"1111111000100111000100",
		b"1111111000100010011011",
		b"1111111000011110000100",
		b"1111111000011001111111",
		b"1111111000010110001011",
		b"1111111000010010101010",
		b"1111111000001111011011",
		b"1111111000001100011111",
		b"1111111000001001110100",
		b"1111111000000111011100",
		b"1111111000000101010110",
		b"1111111000000011100011",
		b"1111111000000010000010",
		b"1111111000000000110011",
		b"1111110111111111110111",
		b"1111110111111111001101",
		b"1111110111111110110101",
		b"1111110111111110110000",
		b"1111110111111110111101",
		b"1111110111111111011100",
		b"1111111000000000001101",
		b"1111111000000001010000",
		b"1111111000000010100101",
		b"1111111000000100001100",
		b"1111111000000110000101",
		b"1111111000001000001111",
		b"1111111000001010101011",
		b"1111111000001101011001",
		b"1111111000010000010111",
		b"1111111000010011100110",
		b"1111111000010111000111",
		b"1111111000011010111000",
		b"1111111000011110111001",
		b"1111111000100011001011",
		b"1111111000100111101110",
		b"1111111000101100100000",
		b"1111111000110001100001",
		b"1111111000110110110011",
		b"1111111000111100010011",
		b"1111111001000010000011",
		b"1111111001001000000001",
		b"1111111001001110001110",
		b"1111111001010100101001",
		b"1111111001011011010011",
		b"1111111001100010001010",
		b"1111111001101001001110",
		b"1111111001110000100000",
		b"1111111001110111111110",
		b"1111111001111111101001",
		b"1111111010000111100000",
		b"1111111010001111100011",
		b"1111111010010111110010",
		b"1111111010100000001100",
		b"1111111010101000110001",
		b"1111111010110001100001",
		b"1111111010111010011011",
		b"1111111011000011011110",
		b"1111111011001100101100",
		b"1111111011010110000011",
		b"1111111011011111100010",
		b"1111111011101001001010",
		b"1111111011110010111010",
		b"1111111011111100110010",
		b"1111111100000110110010",
		b"1111111100010000111000",
		b"1111111100011011000101",
		b"1111111100100101011001",
		b"1111111100101111110010",
		b"1111111100111010010001",
		b"1111111101000100110101",
		b"1111111101001111011101",
		b"1111111101011010001010",
		b"1111111101100100111011",
		b"1111111101101111101111",
		b"1111111101111010100111",
		b"1111111110000101100001",
		b"1111111110010000011110",
		b"1111111110011011011100",
		b"1111111110100110011101",
		b"1111111110110001011110",
		b"1111111110111100100000",
		b"1111111111000111100011",
		b"1111111111010010100101",
		b"1111111111011101101000",
		b"1111111111101000101001",
		b"1111111111110011101001",
		b"1111111111111110101000",
		b"0000000000001001100101",
		b"0000000000010100011111",
		b"0000000000011111010111",
		b"0000000000101010001011",
		b"0000000000110100111100",
		b"0000000000111111101001",
		b"0000000001001010010011",
		b"0000000001010100110111",
		b"0000000001011111010111",
		b"0000000001101001110001",
		b"0000000001110100000110",
		b"0000000001111110010100",
		b"0000000010001000011100",
		b"0000000010010010011110",
		b"0000000010011100011001",
		b"0000000010100110001100",
		b"0000000010101111111000",
		b"0000000010111001011011",
		b"0000000011000010110110",
		b"0000000011001100001001",
		b"0000000011010101010011",
		b"0000000011011110010011",
		b"0000000011100111001010",
		b"0000000011101111110111",
		b"0000000011111000011010",
		b"0000000100000000110011",
		b"0000000100001001000001",
		b"0000000100010001000100",
		b"0000000100011000111100",
		b"0000000100100000101001",
		b"0000000100101000001010",
		b"0000000100101111011111",
		b"0000000100110110101000",
		b"0000000100111101100101",
		b"0000000101000100010101",
		b"0000000101001010111001",
		b"0000000101010001001111",
		b"0000000101010111011001",
		b"0000000101011101010101",
		b"0000000101100011000100",
		b"0000000101101000100101",
		b"0000000101101101111000",
		b"0000000101110010111101",
		b"0000000101110111110101",
		b"0000000101111100011110",
		b"0000000110000000111000",
		b"0000000110000101000101",
		b"0000000110001001000010",
		b"0000000110001100110010",
		b"0000000110010000010010",
		b"0000000110010011100011",
		b"0000000110010110100110",
		b"0000000110011001011010",
		b"0000000110011011111110",
		b"0000000110011110010100",
		b"0000000110100000011011",
		b"0000000110100010010010",
		b"0000000110100011111010",
		b"0000000110100101010011",
		b"0000000110100110011101",
		b"0000000110100111011000",
		b"0000000110101000000011",
		b"0000000110101000100000",
		b"0000000110101000101101",
		b"0000000110101000101011",
		b"0000000110101000011010",
		b"0000000110100111111010",
		b"0000000110100111001100",
		b"0000000110100110001110",
		b"0000000110100101000010",
		b"0000000110100011100110",
		b"0000000110100001111101",
		b"0000000110100000000101",
		b"0000000110011101111110",
		b"0000000110011011101001",
		b"0000000110011001000110",
		b"0000000110010110010101",
		b"0000000110010011010110",
		b"0000000110010000001010",
		b"0000000110001100101111",
		b"0000000110001001001000",
		b"0000000110000101010011",
		b"0000000110000001010001",
		b"0000000101111101000010",
		b"0000000101111000100110",
		b"0000000101110011111110",
		b"0000000101101111001010",
		b"0000000101101010001001",
		b"0000000101100100111101",
		b"0000000101011111100101",
		b"0000000101011010000001",
		b"0000000101010100010011",
		b"0000000101001110011001",
		b"0000000101001000010100",
		b"0000000101000010000101",
		b"0000000100111011101100",
		b"0000000100110101001001",
		b"0000000100101110011011",
		b"0000000100100111100101",
		b"0000000100100000100101",
		b"0000000100011001011101",
		b"0000000100010010001011",
		b"0000000100001010110010",
		b"0000000100000011010000",
		b"0000000011111011100110",
		b"0000000011110011110101",
		b"0000000011101011111101",
		b"0000000011100011111110",
		b"0000000011011011111000",
		b"0000000011010011101100",
		b"0000000011001011011011",
		b"0000000011000011000011",
		b"0000000010111010100110",
		b"0000000010110010000100",
		b"0000000010101001011101",
		b"0000000010100000110010",
		b"0000000010011000000011",
		b"0000000010001111010000",
		b"0000000010000110011001",
		b"0000000001111101100000",
		b"0000000001110100100011",
		b"0000000001101011100100",
		b"0000000001100010100011",
		b"0000000001011001100000",
		b"0000000001010000011100",
		b"0000000001000111010111",
		b"0000000000111110010000",
		b"0000000000110101001001",
		b"0000000000101100000010",
		b"0000000000100010111100",
		b"0000000000011001110101",
		b"0000000000010000101111",
		b"0000000000000111101011",
		b"1111111111111110101000",
		b"1111111111110101100110",
		b"1111111111101100100111",
		b"1111111111100011101001",
		b"1111111111011010101111",
		b"1111111111010001111000",
		b"1111111111001001000011",
		b"1111111111000000010011",
		b"1111111110110111100110",
		b"1111111110101110111101",
		b"1111111110100110011001",
		b"1111111110011101111010",
		b"1111111110010101100000",
		b"1111111110001101001011",
		b"1111111110000100111011",
		b"1111111101111100110010",
		b"1111111101110100101111",
		b"1111111101101100110010",
		b"1111111101100100111011",
		b"1111111101011101001100",
		b"1111111101010101100100",
		b"1111111101001110000011",
		b"1111111101000110101010",
		b"1111111100111111011001",
		b"1111111100111000010000",
		b"1111111100110001010000",
		b"1111111100101010011000",
		b"1111111100100011101001",
		b"1111111100011101000011",
		b"1111111100010110100110",
		b"1111111100010000010011",
		b"1111111100001010001001",
		b"1111111100000100001001",
		b"1111111011111110010011",
		b"1111111011111000101000",
		b"1111111011110011000111",
		b"1111111011101101110000",
		b"1111111011101000100100",
		b"1111111011100011100011",
		b"1111111011011110101100",
		b"1111111011011010000001",
		b"1111111011010101100001",
		b"1111111011010001001101",
		b"1111111011001101000100",
		b"1111111011001001000111",
		b"1111111011000101010101",
		b"1111111011000001101111",
		b"1111111010111110010110",
		b"1111111010111011001000",
		b"1111111010111000000110",
		b"1111111010110101010000",
		b"1111111010110010100111",
		b"1111111010110000001010",
		b"1111111010101101111001",
		b"1111111010101011110100",
		b"1111111010101001111100",
		b"1111111010101000010001",
		b"1111111010100110110010",
		b"1111111010100101011111",
		b"1111111010100100011001",
		b"1111111010100011011111",
		b"1111111010100010110010",
		b"1111111010100010010001",
		b"1111111010100001111101",
		b"1111111010100001110101",
		b"1111111010100001111001",
		b"1111111010100010001010",
		b"1111111010100010100111",
		b"1111111010100011010001",
		b"1111111010100100000110",
		b"1111111010100101001000",
		b"1111111010100110010110",
		b"1111111010100111110000",
		b"1111111010101001010101",
		b"1111111010101011000111",
		b"1111111010101101000100",
		b"1111111010101111001101",
		b"1111111010110001100001",
		b"1111111010110100000001",
		b"1111111010110110101100",
		b"1111111010111001100010",
		b"1111111010111100100011",
		b"1111111010111111101111",
		b"1111111011000011000101",
		b"1111111011000110100110",
		b"1111111011001010010010",
		b"1111111011001110001000",
		b"1111111011010010001000",
		b"1111111011010110010001",
		b"1111111011011010100101",
		b"1111111011011111000010",
		b"1111111011100011101000",
		b"1111111011101000011000",
		b"1111111011101101010001",
		b"1111111011110010010010",
		b"1111111011110111011100",
		b"1111111011111100101110",
		b"1111111100000010001001",
		b"1111111100000111101011",
		b"1111111100001101010101",
		b"1111111100010011000111",
		b"1111111100011001000000",
		b"1111111100011111000000",
		b"1111111100100101000110",
		b"1111111100101011010100",
		b"1111111100110001100111",
		b"1111111100111000000001",
		b"1111111100111110100001",
		b"1111111101000101000110",
		b"1111111101001011110000",
		b"1111111101010010100000",
		b"1111111101011001010101",
		b"1111111101100000001110",
		b"1111111101100111001011",
		b"1111111101101110001101",
		b"1111111101110101010010",
		b"1111111101111100011011",
		b"1111111110000011100111",
		b"1111111110001010110110",
		b"1111111110010010001000",
		b"1111111110011001011101",
		b"1111111110100000110100",
		b"1111111110101000001100",
		b"1111111110101111100111",
		b"1111111110110111000010",
		b"1111111110111110011111",
		b"1111111111000101111101",
		b"1111111111001101011100",
		b"1111111111010100111011",
		b"1111111111011100011010",
		b"1111111111100011111001",
		b"1111111111101011010111",
		b"1111111111110010110101",
		b"1111111111111010010010",
		b"0000000000000001101101",
		b"0000000000001001000111",
		b"0000000000010000100000",
		b"0000000000010111110110",
		b"0000000000011111001010",
		b"0000000000100110011100",
		b"0000000000101101101011",
		b"0000000000110100110111",
		b"0000000000111011111111",
		b"0000000001000011000101",
		b"0000000001001010000110",
		b"0000000001010001000100",
		b"0000000001010111111101",
		b"0000000001011110110010",
		b"0000000001100101100011",
		b"0000000001101100001110",
		b"0000000001110010110101",
		b"0000000001111001010110",
		b"0000000001111111110001",
		b"0000000010000110000111",
		b"0000000010001100010111",
		b"0000000010010010100001",
		b"0000000010011000100100",
		b"0000000010011110100001",
		b"0000000010100100011000",
		b"0000000010101010000111",
		b"0000000010101111101111",
		b"0000000010110101010000",
		b"0000000010111010101010",
		b"0000000010111111111100",
		b"0000000011000101000110",
		b"0000000011001010001000",
		b"0000000011001111000010",
		b"0000000011010011110100",
		b"0000000011011000011110",
		b"0000000011011100111111",
		b"0000000011100001010111",
		b"0000000011100101100111",
		b"0000000011101001101101",
		b"0000000011101101101011",
		b"0000000011110001100000",
		b"0000000011110101001011",
		b"0000000011111000101101",
		b"0000000011111100000101",
		b"0000000011111111010100",
		b"0000000100000010011010",
		b"0000000100000101010110",
		b"0000000100001000001000",
		b"0000000100001010110000",
		b"0000000100001101001110",
		b"0000000100001111100010",
		b"0000000100010001101100",
		b"0000000100010011101101",
		b"0000000100010101100011",
		b"0000000100010111001111",
		b"0000000100011000110001",
		b"0000000100011010001000",
		b"0000000100011011010110",
		b"0000000100011100011001",
		b"0000000100011101010010",
		b"0000000100011110000001",
		b"0000000100011110100101",
		b"0000000100011111000000",
		b"0000000100011111010000",
		b"0000000100011111010110",
		b"0000000100011111010010",
		b"0000000100011111000100",
		b"0000000100011110101011",
		b"0000000100011110001001",
		b"0000000100011101011101",
		b"0000000100011100100111",
		b"0000000100011011100111",
		b"0000000100011010011101",
		b"0000000100011001001001",
		b"0000000100010111101100",
		b"0000000100010110000101",
		b"0000000100010100010101",
		b"0000000100010010011100",
		b"0000000100010000011001",
		b"0000000100001110001101",
		b"0000000100001011110111",
		b"0000000100001001011001",
		b"0000000100000110110010",
		b"0000000100000100000010",
		b"0000000100000001001010",
		b"0000000011111110001001",
		b"0000000011111011000000",
		b"0000000011110111101110",
		b"0000000011110100010101",
		b"0000000011110000110011",
		b"0000000011101101001010",
		b"0000000011101001011001",
		b"0000000011100101100001",
		b"0000000011100001100001",
		b"0000000011011101011010",
		b"0000000011011001001100",
		b"0000000011010100110111",
		b"0000000011010000011100",
		b"0000000011001011111010",
		b"0000000011000111010010",
		b"0000000011000010100100",
		b"0000000010111101110000",
		b"0000000010111000110110",
		b"0000000010110011110110",
		b"0000000010101110110001",
		b"0000000010101001100111",
		b"0000000010100100011000",
		b"0000000010011111000100",
		b"0000000010011001101100",
		b"0000000010010100001111",
		b"0000000010001110101111",
		b"0000000010001001001010",
		b"0000000010000011100001",
		b"0000000001111101110101",
		b"0000000001111000000110",
		b"0000000001110010010011",
		b"0000000001101100011110",
		b"0000000001100110100110",
		b"0000000001100000101011",
		b"0000000001011010101110",
		b"0000000001010100110000",
		b"0000000001001110101111",
		b"0000000001001000101101",
		b"0000000001000010101001",
		b"0000000000111100100100",
		b"0000000000110110011110",
		b"0000000000110000011000",
		b"0000000000101010010001",
		b"0000000000100100001010",
		b"0000000000011110000010",
		b"0000000000010111111011",
		b"0000000000010001110100",
		b"0000000000001011101110",
		b"0000000000000101101000",
		b"1111111111111111100100",
		b"1111111111111001100000",
		b"1111111111110011011110",
		b"1111111111101101011110",
		b"1111111111100111011111",
		b"1111111111100001100011",
		b"1111111111011011101001",
		b"1111111111010101110001",
		b"1111111111001111111100",
		b"1111111111001010001001",
		b"1111111111000100011010",
		b"1111111110111110101110",
		b"1111111110111001000101",
		b"1111111110110011100000",
		b"1111111110101101111110",
		b"1111111110101000100001",
		b"1111111110100011001000",
		b"1111111110011101110011",
		b"1111111110011000100010",
		b"1111111110010011010110",
		b"1111111110001110001111",
		b"1111111110001001001101",
		b"1111111110000100010000",
		b"1111111101111111011001",
		b"1111111101111010100111",
		b"1111111101110101111010",
		b"1111111101110001010100",
		b"1111111101101100110011",
		b"1111111101101000011000",
		b"1111111101100100000100",
		b"1111111101011111110110",
		b"1111111101011011101110",
		b"1111111101010111101101",
		b"1111111101010011110010",
		b"1111111101001111111110",
		b"1111111101001100010010",
		b"1111111101001000101100",
		b"1111111101000101001101",
		b"1111111101000001110110",
		b"1111111100111110100110",
		b"1111111100111011011110",
		b"1111111100111000011101",
		b"1111111100110101100011",
		b"1111111100110010110001",
		b"1111111100110000000111",
		b"1111111100101101100101",
		b"1111111100101011001011",
		b"1111111100101000111000",
		b"1111111100100110101110",
		b"1111111100100100101100",
		b"1111111100100010110001",
		b"1111111100100000111111",
		b"1111111100011111010101",
		b"1111111100011101110100",
		b"1111111100011100011010",
		b"1111111100011011001001",
		b"1111111100011010000000",
		b"1111111100011000111111",
		b"1111111100011000000111",
		b"1111111100010111010111",
		b"1111111100010110101111",
		b"1111111100010110010000",
		b"1111111100010101111001",
		b"1111111100010101101010",
		b"1111111100010101100011",
		b"1111111100010101100101",
		b"1111111100010101101111",
		b"1111111100010110000001",
		b"1111111100010110011011",
		b"1111111100010110111101",
		b"1111111100010111101000",
		b"1111111100011000011010",
		b"1111111100011001010101",
		b"1111111100011010010111",
		b"1111111100011011100001",
		b"1111111100011100110011",
		b"1111111100011110001100",
		b"1111111100011111101110",
		b"1111111100100001010111",
		b"1111111100100011000111",
		b"1111111100100100111111",
		b"1111111100100110111110",
		b"1111111100101001000100",
		b"1111111100101011010001",
		b"1111111100101101100101",
		b"1111111100110000000001",
		b"1111111100110010100011",
		b"1111111100110101001100",
		b"1111111100110111111011",
		b"1111111100111010110001",
		b"1111111100111101101101",
		b"1111111101000000101111",
		b"1111111101000011111000",
		b"1111111101000111000110",
		b"1111111101001010011011",
		b"1111111101001101110101",
		b"1111111101010001010100",
		b"1111111101010100111001",
		b"1111111101011000100011",
		b"1111111101011100010011",
		b"1111111101100000000111",
		b"1111111101100100000001",
		b"1111111101100111111111",
		b"1111111101101100000001",
		b"1111111101110000001000",
		b"1111111101110100010011",
		b"1111111101111000100010",
		b"1111111101111100110101",
		b"1111111110000001001100",
		b"1111111110000101100110",
		b"1111111110001010000100",
		b"1111111110001110100101",
		b"1111111110010011001001",
		b"1111111110010111110000",
		b"1111111110011100011010",
		b"1111111110100001000110",
		b"1111111110100101110100",
		b"1111111110101010100101",
		b"1111111110101111011000",
		b"1111111110110100001101",
		b"1111111110111001000011",
		b"1111111110111101111011",
		b"1111111111000010110101",
		b"1111111111000111101111",
		b"1111111111001100101010",
		b"1111111111010001100111",
		b"1111111111010110100011",
		b"1111111111011011100001",
		b"1111111111100000011110",
		b"1111111111100101011100",
		b"1111111111101010011010",
		b"1111111111101111010111",
		b"1111111111110100010100",
		b"1111111111111001010001",
		b"1111111111111110001100",
		b"0000000000000011000111",
		b"0000000000001000000001",
		b"0000000000001100111001",
		b"0000000000010001110000",
		b"0000000000010110100101",
		b"0000000000011011011001",
		b"0000000000100000001010",
		b"0000000000100100111010",
		b"0000000000101001100111",
		b"0000000000101110010010",
		b"0000000000110010111010",
		b"0000000000110111100000",
		b"0000000000111100000011",
		b"0000000001000000100011",
		b"0000000001000100111111",
		b"0000000001001001011000",
		b"0000000001001101101110",
		b"0000000001010010000000",
		b"0000000001010110001111",
		b"0000000001011010011010",
		b"0000000001011110100000",
		b"0000000001100010100011",
		b"0000000001100110100001",
		b"0000000001101010011011",
		b"0000000001101110010000",
		b"0000000001110010000001",
		b"0000000001110101101101",
		b"0000000001111001010100",
		b"0000000001111100110110",
		b"0000000010000000010011",
		b"0000000010000011101011",
		b"0000000010000110111101",
		b"0000000010001010001010",
		b"0000000010001101010010",
		b"0000000010010000010100",
		b"0000000010010011010001",
		b"0000000010010110000111",
		b"0000000010011000111000",
		b"0000000010011011100011",
		b"0000000010011110001000",
		b"0000000010100000100111",
		b"0000000010100011000000",
		b"0000000010100101010011",
		b"0000000010100111011111",
		b"0000000010101001100101",
		b"0000000010101011100101",
		b"0000000010101101011110",
		b"0000000010101111010001",
		b"0000000010110000111101",
		b"0000000010110010100011",
		b"0000000010110100000011",
		b"0000000010110101011011",
		b"0000000010110110101101",
		b"0000000010110111111001",
		b"0000000010111000111110",
		b"0000000010111001111100",
		b"0000000010111010110011",
		b"0000000010111011100100",
		b"0000000010111100001110",
		b"0000000010111100110001",
		b"0000000010111101001110",
		b"0000000010111101100100",
		b"0000000010111101110011",
		b"0000000010111101111011",
		b"0000000010111101111101",
		b"0000000010111101111001",
		b"0000000010111101101101",
		b"0000000010111101011011",
		b"0000000010111101000011",
		b"0000000010111100100100",
		b"0000000010111011111110",
		b"0000000010111011010010",
		b"0000000010111010100000",
		b"0000000010111001100111",
		b"0000000010111000101000",
		b"0000000010110111100010",
		b"0000000010110110010111",
		b"0000000010110101000101",
		b"0000000010110011101110",
		b"0000000010110010010000",
		b"0000000010110000101100",
		b"0000000010101111000011",
		b"0000000010101101010100",
		b"0000000010101011011111",
		b"0000000010101001100100",
		b"0000000010100111100100",
		b"0000000010100101011111",
		b"0000000010100011010100",
		b"0000000010100001000100",
		b"0000000010011110101111",
		b"0000000010011100010100",
		b"0000000010011001110101",
		b"0000000010010111010001",
		b"0000000010010100101000",
		b"0000000010010001111011",
		b"0000000010001111001001",
		b"0000000010001100010010",
		b"0000000010001001010111",
		b"0000000010000110011000",
		b"0000000010000011010101",
		b"0000000010000000001110",
		b"0000000001111101000011",
		b"0000000001111001110101",
		b"0000000001110110100011",
		b"0000000001110011001101",
		b"0000000001101111110100",
		b"0000000001101100011000",
		b"0000000001101000111001",
		b"0000000001100101010111",
		b"0000000001100001110010",
		b"0000000001011110001010",
		b"0000000001011010100000",
		b"0000000001010110110011",
		b"0000000001010011000101",
		b"0000000001001111010100",
		b"0000000001001011100001",
		b"0000000001000111101100",
		b"0000000001000011110101",
		b"0000000000111111111101",
		b"0000000000111100000100",
		b"0000000000111000001001",
		b"0000000000110100001101",
		b"0000000000110000010000",
		b"0000000000101100010010",
		b"0000000000101000010100",
		b"0000000000100100010101",
		b"0000000000100000010101",
		b"0000000000011100010101",
		b"0000000000011000010101",
		b"0000000000010100010101",
		b"0000000000010000010101",
		b"0000000000001100010101",
		b"0000000000001000010110",
		b"0000000000000100010111",
		b"0000000000000000011001",
		b"1111111111111100011100",
		b"1111111111111000100000",
		b"1111111111110100100101",
		b"1111111111110000101011",
		b"1111111111101100110010",
		b"1111111111101000111011",
		b"1111111111100101000101",
		b"1111111111100001010001",
		b"1111111111011101011111",
		b"1111111111011001101111",
		b"1111111111010110000001",
		b"1111111111010010010110",
		b"1111111111001110101100",
		b"1111111111001011000101",
		b"1111111111000111100001",
		b"1111111111000100000000",
		b"1111111111000000100001",
		b"1111111110111101000101",
		b"1111111110111001101100",
		b"1111111110110110010111",
		b"1111111110110011000100",
		b"1111111110101111110101",
		b"1111111110101100101010",
		b"1111111110101001100010",
		b"1111111110100110011101",
		b"1111111110100011011101",
		b"1111111110100000100000",
		b"1111111110011101100111",
		b"1111111110011010110011",
		b"1111111110011000000010",
		b"1111111110010101010110",
		b"1111111110010010101101",
		b"1111111110010000001010",
		b"1111111110001101101010",
		b"1111111110001011001111",
		b"1111111110001000111001",
		b"1111111110000110100111",
		b"1111111110000100011010",
		b"1111111110000010010010",
		b"1111111110000000001110",
		b"1111111101111110010000",
		b"1111111101111100010110",
		b"1111111101111010100010",
		b"1111111101111000110010",
		b"1111111101110111000111",
		b"1111111101110101100010",
		b"1111111101110100000010",
		b"1111111101110010100110",
		b"1111111101110001010000",
		b"1111111101110000000000",
		b"1111111101101110110100",
		b"1111111101101101101110",
		b"1111111101101100101101",
		b"1111111101101011110010",
		b"1111111101101010111100",
		b"1111111101101010001011",
		b"1111111101101001100000",
		b"1111111101101000111001",
		b"1111111101101000011001",
		b"1111111101100111111110",
		b"1111111101100111101000",
		b"1111111101100111010111",
		b"1111111101100111001100",
		b"1111111101100111000110",
		b"1111111101100111000101",
		b"1111111101100111001010",
		b"1111111101100111010100",
		b"1111111101100111100100",
		b"1111111101100111111000",
		b"1111111101101000010010",
		b"1111111101101000110001",
		b"1111111101101001010101",
		b"1111111101101001111110",
		b"1111111101101010101100",
		b"1111111101101011100000",
		b"1111111101101100011000",
		b"1111111101101101010101",
		b"1111111101101110010111",
		b"1111111101101111011110",
		b"1111111101110000101010",
		b"1111111101110001111011",
		b"1111111101110011010000",
		b"1111111101110100101010",
		b"1111111101110110001000",
		b"1111111101110111101011",
		b"1111111101111001010010",
		b"1111111101111010111101",
		b"1111111101111100101101",
		b"1111111101111110100001",
		b"1111111110000000011001",
		b"1111111110000010010101",
		b"1111111110000100010101",
		b"1111111110000110011001",
		b"1111111110001000100001",
		b"1111111110001010101100",
		b"1111111110001100111011",
		b"1111111110001111001101",
		b"1111111110010001100011",
		b"1111111110010011111100",
		b"1111111110010110011001",
		b"1111111110011000111000",
		b"1111111110011011011011",
		b"1111111110011110000001",
		b"1111111110100000101001",
		b"1111111110100011010100",
		b"1111111110100110000010",
		b"1111111110101000110010",
		b"1111111110101011100101",
		b"1111111110101110011010",
		b"1111111110110001010010",
		b"1111111110110100001011",
		b"1111111110110111000111",
		b"1111111110111010000100",
		b"1111111110111101000011",
		b"1111111111000000000100",
		b"1111111111000011000110",
		b"1111111111000110001010",
		b"1111111111001001001111",
		b"1111111111001100010110",
		b"1111111111001111011101",
		b"1111111111010010100110",
		b"1111111111010101110000",
		b"1111111111011000111010",
		b"1111111111011100000101",
		b"1111111111011111010000",
		b"1111111111100010011100",
		b"1111111111100101101000",
		b"1111111111101000110101",
		b"1111111111101100000010",
		b"1111111111101111001110",
		b"1111111111110010011011",
		b"1111111111110101100111",
		b"1111111111111000110011",
		b"1111111111111011111111",
		b"1111111111111111001010",
		b"0000000000000010010100",
		b"0000000000000101011110",
		b"0000000000001000100110",
		b"0000000000001011101110",
		b"0000000000001110110101",
		b"0000000000010001111010",
		b"0000000000010100111110",
		b"0000000000011000000001",
		b"0000000000011011000010",
		b"0000000000011110000010",
		b"0000000000100001000000",
		b"0000000000100011111100",
		b"0000000000100110110111",
		b"0000000000101001101111",
		b"0000000000101100100101",
		b"0000000000101111011010",
		b"0000000000110010001011",
		b"0000000000110100111011",
		b"0000000000110111101000",
		b"0000000000111010010011",
		b"0000000000111100111011",
		b"0000000000111111100000",
		b"0000000001000010000011",
		b"0000000001000100100010",
		b"0000000001000110111111",
		b"0000000001001001011001",
		b"0000000001001011110000",
		b"0000000001001110000011",
		b"0000000001010000010100",
		b"0000000001010010100001",
		b"0000000001010100101011",
		b"0000000001010110110001",
		b"0000000001011000110100",
		b"0000000001011010110100",
		b"0000000001011100110000",
		b"0000000001011110101000",
		b"0000000001100000011100",
		b"0000000001100010001101",
		b"0000000001100011111010",
		b"0000000001100101100011",
		b"0000000001100111001001",
		b"0000000001101000101010",
		b"0000000001101010001000",
		b"0000000001101011100001",
		b"0000000001101100110110",
		b"0000000001101110001000",
		b"0000000001101111010101",
		b"0000000001110000011110",
		b"0000000001110001100011",
		b"0000000001110010100100",
		b"0000000001110011100001",
		b"0000000001110100011001",
		b"0000000001110101001110",
		b"0000000001110101111110",
		b"0000000001110110101001",
		b"0000000001110111010001",
		b"0000000001110111110100",
		b"0000000001111000010011",
		b"0000000001111000101110",
		b"0000000001111001000100",
		b"0000000001111001010111",
		b"0000000001111001100101",
		b"0000000001111001101110",
		b"0000000001111001110100",
		b"0000000001111001110101",
		b"0000000001111001110010",
		b"0000000001111001101011",
		b"0000000001111001011111",
		b"0000000001111001010000",
		b"0000000001111000111100",
		b"0000000001111000100100",
		b"0000000001111000001000",
		b"0000000001110111101000",
		b"0000000001110111000100",
		b"0000000001110110011100",
		b"0000000001110101110000",
		b"0000000001110101000000",
		b"0000000001110100001101",
		b"0000000001110011010101",
		b"0000000001110010011010",
		b"0000000001110001011010",
		b"0000000001110000011000",
		b"0000000001101111010001",
		b"0000000001101110000111",
		b"0000000001101100111001",
		b"0000000001101011101000",
		b"0000000001101010010100",
		b"0000000001101000111100",
		b"0000000001100111100000",
		b"0000000001100110000010",
		b"0000000001100100100000",
		b"0000000001100010111011",
		b"0000000001100001010011",
		b"0000000001011111101000",
		b"0000000001011101111010",
		b"0000000001011100001001",
		b"0000000001011010010101",
		b"0000000001011000011111",
		b"0000000001010110100110",
		b"0000000001010100101010",
		b"0000000001010010101100",
		b"0000000001010000101100",
		b"0000000001001110101001",
		b"0000000001001100100100",
		b"0000000001001010011101",
		b"0000000001001000010011",
		b"0000000001000110001000",
		b"0000000001000011111010",
		b"0000000001000001101011",
		b"0000000000111111011010",
		b"0000000000111101000111",
		b"0000000000111010110011",
		b"0000000000111000011101",
		b"0000000000110110000110",
		b"0000000000110011101101",
		b"0000000000110001010011",
		b"0000000000101110111000",
		b"0000000000101100011100",
		b"0000000000101001111110",
		b"0000000000100111100000",
		b"0000000000100101000001",
		b"0000000000100010100010",
		b"0000000000100000000001",
		b"0000000000011101100000",
		b"0000000000011010111111",
		b"0000000000011000011101",
		b"0000000000010101111011",
		b"0000000000010011011001",
		b"0000000000010000110111",
		b"0000000000001110010100",
		b"0000000000001011110010",
		b"0000000000001001010000",
		b"0000000000000110101110",
		b"0000000000000100001100",
		b"0000000000000001101011",
		b"1111111111111111001010",
		b"1111111111111100101010",
		b"1111111111111010001011",
		b"1111111111110111101100",
		b"1111111111110101001110",
		b"1111111111110010110001",
		b"1111111111110000010101",
		b"1111111111101101111010",
		b"1111111111101011100000",
		b"1111111111101001001000",
		b"1111111111100110110000",
		b"1111111111100100011010",
		b"1111111111100010000110",
		b"1111111111011111110011",
		b"1111111111011101100010",
		b"1111111111011011010010",
		b"1111111111011001000100",
		b"1111111111010110111000",
		b"1111111111010100101110",
		b"1111111111010010100110",
		b"1111111111010000100000",
		b"1111111111001110011100",
		b"1111111111001100011010",
		b"1111111111001010011010",
		b"1111111111001000011100",
		b"1111111111000110100001",
		b"1111111111000100101001",
		b"1111111111000010110010",
		b"1111111111000000111111",
		b"1111111110111111001101",
		b"1111111110111101011111",
		b"1111111110111011110011",
		b"1111111110111010001010",
		b"1111111110111000100011",
		b"1111111110110110111111",
		b"1111111110110101011111",
		b"1111111110110100000001",
		b"1111111110110010100110",
		b"1111111110110001001110",
		b"1111111110101111111001",
		b"1111111110101110100111",
		b"1111111110101101011000",
		b"1111111110101100001100",
		b"1111111110101011000011",
		b"1111111110101001111110",
		b"1111111110101000111011",
		b"1111111110100111111100",
		b"1111111110100111000000",
		b"1111111110100110000111",
		b"1111111110100101010010",
		b"1111111110100100100000",
		b"1111111110100011110001",
		b"1111111110100011000110",
		b"1111111110100010011110",
		b"1111111110100001111001",
		b"1111111110100001010111",
		b"1111111110100000111001",
		b"1111111110100000011110",
		b"1111111110100000000111",
		b"1111111110011111110011",
		b"1111111110011111100010",
		b"1111111110011111010101",
		b"1111111110011111001011",
		b"1111111110011111000100",
		b"1111111110011111000001",
		b"1111111110011111000001",
		b"1111111110011111000100",
		b"1111111110011111001011",
		b"1111111110011111010101",
		b"1111111110011111100010",
		b"1111111110011111110011",
		b"1111111110100000000110",
		b"1111111110100000011101",
		b"1111111110100000110111",
		b"1111111110100001010101",
		b"1111111110100001110101",
		b"1111111110100010011000",
		b"1111111110100010111111",
		b"1111111110100011101000",
		b"1111111110100100010101",
		b"1111111110100101000101",
		b"1111111110100101110111",
		b"1111111110100110101100",
		b"1111111110100111100101",
		b"1111111110101000100000",
		b"1111111110101001011110",
		b"1111111110101010011110",
		b"1111111110101011100001",
		b"1111111110101100100111",
		b"1111111110101101110000",
		b"1111111110101110111011",
		b"1111111110110000001000",
		b"1111111110110001011000",
		b"1111111110110010101011",
		b"1111111110110100000000",
		b"1111111110110101010111",
		b"1111111110110110110000",
		b"1111111110111000001011",
		b"1111111110111001101001",
		b"1111111110111011001001",
		b"1111111110111100101010",
		b"1111111110111110001110",
		b"1111111110111111110011",
		b"1111111111000001011011",
		b"1111111111000011000100",
		b"1111111111000100101110",
		b"1111111111000110011011",
		b"1111111111001000001001",
		b"1111111111001001111000",
		b"1111111111001011101001",
		b"1111111111001101011011",
		b"1111111111001111001111",
		b"1111111111010001000100",
		b"1111111111010010111010",
		b"1111111111010100110001",
		b"1111111111010110101001",
		b"1111111111011000100010",
		b"1111111111011010011100",
		b"1111111111011100010111",
		b"1111111111011110010011",
		b"1111111111100000001111",
		b"1111111111100010001100",
		b"1111111111100100001010",
		b"1111111111100110001000",
		b"1111111111101000000111",
		b"1111111111101010000101",
		b"1111111111101100000100",
		b"1111111111101110000100",
		b"1111111111110000000011",
		b"1111111111110010000011",
		b"1111111111110100000010",
		b"1111111111110110000010",
		b"1111111111111000000001",
		b"1111111111111010000000",
		b"1111111111111011111111",
		b"1111111111111101111110",
		b"1111111111111111111100",
		b"0000000000000001111010",
		b"0000000000000011110111",
		b"0000000000000101110100",
		b"0000000000000111110000",
		b"0000000000001001101011",
		b"0000000000001011100101",
		b"0000000000001101011111",
		b"0000000000001111011000",
		b"0000000000010001001111",
		b"0000000000010011000110",
		b"0000000000010100111100",
		b"0000000000010110110000",
		b"0000000000011000100011",
		b"0000000000011010010101",
		b"0000000000011100000110",
		b"0000000000011101110101",
		b"0000000000011111100011",
		b"0000000000100001001111",
		b"0000000000100010111010",
		b"0000000000100100100011",
		b"0000000000100110001011",
		b"0000000000100111110001",
		b"0000000000101001010101",
		b"0000000000101010110111",
		b"0000000000101100011000",
		b"0000000000101101110111",
		b"0000000000101111010011",
		b"0000000000110000101110",
		b"0000000000110010000111",
		b"0000000000110011011110",
		b"0000000000110100110010",
		b"0000000000110110000101",
		b"0000000000110111010101",
		b"0000000000111000100011",
		b"0000000000111001101111",
		b"0000000000111010111001",
		b"0000000000111100000000",
		b"0000000000111101000101",
		b"0000000000111110001000",
		b"0000000000111111001001",
		b"0000000001000000000111",
		b"0000000001000001000010",
		b"0000000001000001111011",
		b"0000000001000010110010",
		b"0000000001000011100110",
		b"0000000001000100010111",
		b"0000000001000101000111",
		b"0000000001000101110011",
		b"0000000001000110011101",
		b"0000000001000111000100",
		b"0000000001000111101001",
		b"0000000001001000001100",
		b"0000000001001000101011",
		b"0000000001001001001000",
		b"0000000001001001100011",
		b"0000000001001001111010",
		b"0000000001001010001111",
		b"0000000001001010100010",
		b"0000000001001010110010",
		b"0000000001001010111111",
		b"0000000001001011001010",
		b"0000000001001011010010",
		b"0000000001001011010111",
		b"0000000001001011011010",
		b"0000000001001011011010",
		b"0000000001001011011000",
		b"0000000001001011010011",
		b"0000000001001011001011",
		b"0000000001001011000001",
		b"0000000001001010110101",
		b"0000000001001010100110",
		b"0000000001001010010100",
		b"0000000001001010000000",
		b"0000000001001001101001",
		b"0000000001001001010000",
		b"0000000001001000110101",
		b"0000000001001000010111",
		b"0000000001000111110110",
		b"0000000001000111010100",
		b"0000000001000110101111",
		b"0000000001000110001000",
		b"0000000001000101011110",
		b"0000000001000100110010",
		b"0000000001000100000100",
		b"0000000001000011010100",
		b"0000000001000010100010",
		b"0000000001000001101101",
		b"0000000001000000110111",
		b"0000000000111111111111",
		b"0000000000111111000100",
		b"0000000000111110001000",
		b"0000000000111101001001",
		b"0000000000111100001001",
		b"0000000000111011000111",
		b"0000000000111010000011",
		b"0000000000111000111101",
		b"0000000000110111110110",
		b"0000000000110110101101",
		b"0000000000110101100010",
		b"0000000000110100010110",
		b"0000000000110011001000",
		b"0000000000110001111001",
		b"0000000000110000101000",
		b"0000000000101111010110",
		b"0000000000101110000010",
		b"0000000000101100101110",
		b"0000000000101011011000",
		b"0000000000101010000001",
		b"0000000000101000101000",
		b"0000000000100111001111",
		b"0000000000100101110100",
		b"0000000000100100011001",
		b"0000000000100010111100",
		b"0000000000100001011111",
		b"0000000000100000000001",
		b"0000000000011110100010",
		b"0000000000011101000011",
		b"0000000000011011100010",
		b"0000000000011010000001",
		b"0000000000011000100000",
		b"0000000000010110111110",
		b"0000000000010101011011",
		b"0000000000010011111001",
		b"0000000000010010010101",
		b"0000000000010000110010",
		b"0000000000001111001110",
		b"0000000000001101101010",
		b"0000000000001100000110",
		b"0000000000001010100010",
		b"0000000000001000111101",
		b"0000000000000111011001",
		b"0000000000000101110101",
		b"0000000000000100010001",
		b"0000000000000010101101",
		b"0000000000000001001010",
		b"1111111111111111100110",
		b"1111111111111110000011",
		b"1111111111111100100001",
		b"1111111111111010111111",
		b"1111111111111001011101",
		b"1111111111110111111100",
		b"1111111111110110011011",
		b"1111111111110100111011",
		b"1111111111110011011100",
		b"1111111111110001111101",
		b"1111111111110000100000",
		b"1111111111101111000011",
		b"1111111111101101100111",
		b"1111111111101100001100",
		b"1111111111101010110001",
		b"1111111111101001011000",
		b"1111111111101000000000",
		b"1111111111100110101001",
		b"1111111111100101010011",
		b"1111111111100011111110",
		b"1111111111100010101011",
		b"1111111111100001011000",
		b"1111111111100000000111",
		b"1111111111011110111000",
		b"1111111111011101101001",
		b"1111111111011100011100",
		b"1111111111011011010001",
		b"1111111111011010000111",
		b"1111111111011000111110",
		b"1111111111010111110111",
		b"1111111111010110110010",
		b"1111111111010101101110",
		b"1111111111010100101100",
		b"1111111111010011101100",
		b"1111111111010010101101",
		b"1111111111010001110000",
		b"1111111111010000110100",
		b"1111111111001111111011",
		b"1111111111001111000011",
		b"1111111111001110001101",
		b"1111111111001101011000",
		b"1111111111001100100110",
		b"1111111111001011110110",
		b"1111111111001011000111",
		b"1111111111001010011010",
		b"1111111111001001110000",
		b"1111111111001001000111",
		b"1111111111001000100000",
		b"1111111111000111111011",
		b"1111111111000111011000",
		b"1111111111000110110111",
		b"1111111111000110011000",
		b"1111111111000101111011",
		b"1111111111000101100000",
		b"1111111111000101000111",
		b"1111111111000100110000",
		b"1111111111000100011100",
		b"1111111111000100001001",
		b"1111111111000011111000",
		b"1111111111000011101001",
		b"1111111111000011011101",
		b"1111111111000011010010",
		b"1111111111000011001001",
		b"1111111111000011000011",
		b"1111111111000010111110",
		b"1111111111000010111100",
		b"1111111111000010111011",
		b"1111111111000010111101",
		b"1111111111000011000000",
		b"1111111111000011000101",
		b"1111111111000011001101",
		b"1111111111000011010110",
		b"1111111111000011100010",
		b"1111111111000011101111",
		b"1111111111000011111110",
		b"1111111111000100010000",
		b"1111111111000100100011",
		b"1111111111000100111000",
		b"1111111111000101001110",
		b"1111111111000101100111",
		b"1111111111000110000010",
		b"1111111111000110011110",
		b"1111111111000110111100",
		b"1111111111000111011100",
		b"1111111111000111111101",
		b"1111111111001000100001",
		b"1111111111001001000110",
		b"1111111111001001101100",
		b"1111111111001010010100",
		b"1111111111001010111110",
		b"1111111111001011101010",
		b"1111111111001100010111",
		b"1111111111001101000101",
		b"1111111111001101110101",
		b"1111111111001110100111",
		b"1111111111001111011010",
		b"1111111111010000001110",
		b"1111111111010001000100",
		b"1111111111010001111011",
		b"1111111111010010110011",
		b"1111111111010011101101",
		b"1111111111010100100111",
		b"1111111111010101100011",
		b"1111111111010110100001",
		b"1111111111010111011111",
		b"1111111111011000011110",
		b"1111111111011001011111",
		b"1111111111011010100000",
		b"1111111111011011100010",
		b"1111111111011100100110",
		b"1111111111011101101010",
		b"1111111111011110101111",
		b"1111111111011111110101",
		b"1111111111100000111011",
		b"1111111111100010000011",
		b"1111111111100011001011",
		b"1111111111100100010011",
		b"1111111111100101011101",
		b"1111111111100110100111",
		b"1111111111100111110001",
		b"1111111111101000111100",
		b"1111111111101010000111",
		b"1111111111101011010011",
		b"1111111111101100011111",
		b"1111111111101101101100",
		b"1111111111101110111000",
		b"1111111111110000000101",
		b"1111111111110001010011",
		b"1111111111110010100000",
		b"1111111111110011101101",
		b"1111111111110100111011",
		b"1111111111110110001000",
		b"1111111111110111010110",
		b"1111111111111000100100",
		b"1111111111111001110001",
		b"1111111111111010111110",
		b"1111111111111100001011",
		b"1111111111111101011000",
		b"1111111111111110100101",
		b"1111111111111111110001",
		b"0000000000000000111101",
		b"0000000000000010001001",
		b"0000000000000011010100",
		b"0000000000000100011111",
		b"0000000000000101101010",
		b"0000000000000110110100",
		b"0000000000000111111101",
		b"0000000000001001000110",
		b"0000000000001010001110",
		b"0000000000001011010101",
		b"0000000000001100011100",
		b"0000000000001101100010",
		b"0000000000001110100111",
		b"0000000000001111101011",
		b"0000000000010000101111",
		b"0000000000010001110010",
		b"0000000000010010110100",
		b"0000000000010011110101",
		b"0000000000010100110100",
		b"0000000000010101110011",
		b"0000000000010110110001",
		b"0000000000010111101110",
		b"0000000000011000101010",
		b"0000000000011001100101",
		b"0000000000011010011110",
		b"0000000000011011010111",
		b"0000000000011100001110",
		b"0000000000011101000100",
		b"0000000000011101111001",
		b"0000000000011110101100",
		b"0000000000011111011111",
		b"0000000000100000010000",
		b"0000000000100000111111",
		b"0000000000100001101101",
		b"0000000000100010011010",
		b"0000000000100011000110",
		b"0000000000100011110000",
		b"0000000000100100011001",
		b"0000000000100101000000",
		b"0000000000100101100110",
		b"0000000000100110001010",
		b"0000000000100110101101",
		b"0000000000100111001111",
		b"0000000000100111101111",
		b"0000000000101000001101",
		b"0000000000101000101010",
		b"0000000000101001000101",
		b"0000000000101001011111",
		b"0000000000101001110111",
		b"0000000000101010001110",
		b"0000000000101010100011",
		b"0000000000101010110110",
		b"0000000000101011001000",
		b"0000000000101011011001",
		b"0000000000101011101000",
		b"0000000000101011110101",
		b"0000000000101100000000",
		b"0000000000101100001010",
		b"0000000000101100010011",
		b"0000000000101100011001",
		b"0000000000101100011111",
		b"0000000000101100100010",
		b"0000000000101100100100",
		b"0000000000101100100101",
		b"0000000000101100100100",
		b"0000000000101100100001",
		b"0000000000101100011101",
		b"0000000000101100010111",
		b"0000000000101100010000",
		b"0000000000101100000111",
		b"0000000000101011111100",
		b"0000000000101011110000",
		b"0000000000101011100011",
		b"0000000000101011010100",
		b"0000000000101011000011",
		b"0000000000101010110001",
		b"0000000000101010011110",
		b"0000000000101010001001",
		b"0000000000101001110011",
		b"0000000000101001011011",
		b"0000000000101001000010",
		b"0000000000101000101000",
		b"0000000000101000001100",
		b"0000000000100111101111",
		b"0000000000100111010000",
		b"0000000000100110110000",
		b"0000000000100110001111",
		b"0000000000100101101101",
		b"0000000000100101001001",
		b"0000000000100100100101",
		b"0000000000100011111110",
		b"0000000000100011010111",
		b"0000000000100010101111",
		b"0000000000100010000101",
		b"0000000000100001011011",
		b"0000000000100000101111",
		b"0000000000100000000010",
		b"0000000000011111010101",
		b"0000000000011110100110",
		b"0000000000011101110110",
		b"0000000000011101000101",
		b"0000000000011100010100",
		b"0000000000011011100001",
		b"0000000000011010101110",
		b"0000000000011001111010",
		b"0000000000011001000101",
		b"0000000000011000001111",
		b"0000000000010111011000",
		b"0000000000010110100001",
		b"0000000000010101101001",
		b"0000000000010100110001",
		b"0000000000010011110111",
		b"0000000000010010111110",
		b"0000000000010010000011",
		b"0000000000010001001000",
		b"0000000000010000001101",
		b"0000000000001111010001",
		b"0000000000001110010101",
		b"0000000000001101011000",
		b"0000000000001100011011",
		b"0000000000001011011101",
		b"0000000000001010011111",
		b"0000000000001001100001",
		b"0000000000001000100011",
		b"0000000000000111100100",
		b"0000000000000110100110",
		b"0000000000000101100111",
		b"0000000000000100101000",
		b"0000000000000011101001",
		b"0000000000000010101001",
		b"0000000000000001101010",
		b"0000000000000000101011",
		b"1111111111111111101100",
		b"1111111111111110101101",
		b"1111111111111101101110",
		b"1111111111111100101111",
		b"1111111111111011110000",
		b"1111111111111010110010",
		b"1111111111111001110011",
		b"1111111111111000110101",
		b"1111111111110111110111",
		b"1111111111110110111010",
		b"1111111111110101111101",
		b"1111111111110101000000",
		b"1111111111110100000100",
		b"1111111111110011001000",
		b"1111111111110010001100",
		b"1111111111110001010001",
		b"1111111111110000010111",
		b"1111111111101111011101",
		b"1111111111101110100100",
		b"1111111111101101101011",
		b"1111111111101100110011",
		b"1111111111101011111011",
		b"1111111111101011000100",
		b"1111111111101010001110",
		b"1111111111101001011001",
		b"1111111111101000100100",
		b"1111111111100111110000",
		b"1111111111100110111101",
		b"1111111111100110001010",
		b"1111111111100101011001",
		b"1111111111100100101000",
		b"1111111111100011111000",
		b"1111111111100011001001",
		b"1111111111100010011011",
		b"1111111111100001101110",
		b"1111111111100001000010",
		b"1111111111100000010111",
		b"1111111111011111101101",
		b"1111111111011111000100",
		b"1111111111011110011100",
		b"1111111111011101110101",
		b"1111111111011101001111",
		b"1111111111011100101010",
		b"1111111111011100000110",
		b"1111111111011011100011",
		b"1111111111011011000010",
		b"1111111111011010100001",
		b"1111111111011010000010",
		b"1111111111011001100100",
		b"1111111111011001000110",
		b"1111111111011000101011",
		b"1111111111011000010000",
		b"1111111111010111110110",
		b"1111111111010111011110",
		b"1111111111010111000111",
		b"1111111111010110110001",
		b"1111111111010110011100",
		b"1111111111010110001001",
		b"1111111111010101110111",
		b"1111111111010101100110",
		b"1111111111010101010110",
		b"1111111111010101000111",
		b"1111111111010100111010",
		b"1111111111010100101110",
		b"1111111111010100100011",
		b"1111111111010100011010",
		b"1111111111010100010001",
		b"1111111111010100001010",
		b"1111111111010100000101",
		b"1111111111010100000000",
		b"1111111111010011111101",
		b"1111111111010011111011",
		b"1111111111010011111010",
		b"1111111111010011111010",
		b"1111111111010011111100",
		b"1111111111010011111111",
		b"1111111111010100000011",
		b"1111111111010100001000",
		b"1111111111010100001110",
		b"1111111111010100010110",
		b"1111111111010100011111",
		b"1111111111010100101001",
		b"1111111111010100110100",
		b"1111111111010101000001",
		b"1111111111010101001110",
		b"1111111111010101011101",
		b"1111111111010101101101",
		b"1111111111010101111101",
		b"1111111111010110001111",
		b"1111111111010110100011",
		b"1111111111010110110111",
		b"1111111111010111001100",
		b"1111111111010111100010",
		b"1111111111010111111010",
		b"1111111111011000010010",
		b"1111111111011000101011",
		b"1111111111011001000101",
		b"1111111111011001100001",
		b"1111111111011001111101",
		b"1111111111011010011010",
		b"1111111111011010111000",
		b"1111111111011011010111",
		b"1111111111011011110111",
		b"1111111111011100011000",
		b"1111111111011100111001",
		b"1111111111011101011100",
		b"1111111111011101111111",
		b"1111111111011110100011",
		b"1111111111011111001000",
		b"1111111111011111101101",
		b"1111111111100000010011",
		b"1111111111100000111010",
		b"1111111111100001100010",
		b"1111111111100010001010",
		b"1111111111100010110011",
		b"1111111111100011011100",
		b"1111111111100100000110",
		b"1111111111100100110001",
		b"1111111111100101011100",
		b"1111111111100110000111",
		b"1111111111100110110011",
		b"1111111111100111100000",
		b"1111111111101000001101",
		b"1111111111101000111010",
		b"1111111111101001101000",
		b"1111111111101010010110",
		b"1111111111101011000101",
		b"1111111111101011110100",
		b"1111111111101100100011",
		b"1111111111101101010010",
		b"1111111111101110000010",
		b"1111111111101110110010",
		b"1111111111101111100010",
		b"1111111111110000010010",
		b"1111111111110001000011",
		b"1111111111110001110011",
		b"1111111111110010100100",
		b"1111111111110011010100",
		b"1111111111110100000101",
		b"1111111111110100110110",
		b"1111111111110101100111",
		b"1111111111110110010111",
		b"1111111111110111001000",
		b"1111111111110111111001",
		b"1111111111111000101001",
		b"1111111111111001011010",
		b"1111111111111010001010",
		b"1111111111111010111010",
		b"1111111111111011101010",
		b"1111111111111100011001",
		b"1111111111111101001001",
		b"1111111111111101111000",
		b"1111111111111110100111",
		b"1111111111111111010101",
		b"0000000000000000000011",
		b"0000000000000000110001",
		b"0000000000000001011110",
		b"0000000000000010001011",
		b"0000000000000010111000",
		b"0000000000000011100100",
		b"0000000000000100010000",
		b"0000000000000100111011",
		b"0000000000000101100110",
		b"0000000000000110010000",
		b"0000000000000110111001",
		b"0000000000000111100011",
		b"0000000000001000001011",
		b"0000000000001000110011",
		b"0000000000001001011010",
		b"0000000000001010000000",
		b"0000000000001010100110",
		b"0000000000001011001100",
		b"0000000000001011110000",
		b"0000000000001100010100",
		b"0000000000001100110111",
		b"0000000000001101011001",
		b"0000000000001101111011",
		b"0000000000001110011011",
		b"0000000000001110111011",
		b"0000000000001111011010",
		b"0000000000001111111001",
		b"0000000000010000010110",
		b"0000000000010000110011",
		b"0000000000010001001111",
		b"0000000000010001101001",
		b"0000000000010010000011",
		b"0000000000010010011100",
		b"0000000000010010110101",
		b"0000000000010011001100",
		b"0000000000010011100010",
		b"0000000000010011110111",
		b"0000000000010100001100",
		b"0000000000010100011111",
		b"0000000000010100110010",
		b"0000000000010101000011",
		b"0000000000010101010100",
		b"0000000000010101100011",
		b"0000000000010101110010",
		b"0000000000010101111111",
		b"0000000000010110001011",
		b"0000000000010110010111",
		b"0000000000010110100001",
		b"0000000000010110101011",
		b"0000000000010110110011",
		b"0000000000010110111010",
		b"0000000000010111000000",
		b"0000000000010111000110",
		b"0000000000010111001010",
		b"0000000000010111001101",
		b"0000000000010111001111",
		b"0000000000010111010000",
		b"0000000000010111010000",
		b"0000000000010111001111",
		b"0000000000010111001100",
		b"0000000000010111001001",
		b"0000000000010111000101",
		b"0000000000010111000000",
		b"0000000000010110111001",
		b"0000000000010110110010",
		b"0000000000010110101001",
		b"0000000000010110100000",
		b"0000000000010110010110",
		b"0000000000010110001010",
		b"0000000000010101111101",
		b"0000000000010101110000",
		b"0000000000010101100001",
		b"0000000000010101010010",
		b"0000000000010101000001",
		b"0000000000010100110000",
		b"0000000000010100011101",
		b"0000000000010100001010",
		b"0000000000010011110101",
		b"0000000000010011100000",
		b"0000000000010011001001",
		b"0000000000010010110010",
		b"0000000000010010011010",
		b"0000000000010010000001",
		b"0000000000010001100111",
		b"0000000000010001001100",
		b"0000000000010000110000",
		b"0000000000010000010011",
		b"0000000000001111110110",
		b"0000000000001111010111",
		b"0000000000001110111000",
		b"0000000000001110011000",
		b"0000000000001101110111",
		b"0000000000001101010101",
		b"0000000000001100110011",
		b"0000000000001100001111",
		b"0000000000001011101011",
		b"0000000000001011000111",
		b"0000000000001010100001",
		b"0000000000001001111011",
		b"0000000000001001010100",
		b"0000000000001000101101",
		b"0000000000001000000101",
		b"0000000000000111011100",
		b"0000000000000110110010",
		b"0000000000000110001000",
		b"0000000000000101011101",
		b"0000000000000100110010",
		b"0000000000000100000110",
		b"0000000000000011011010",
		b"0000000000000010101101",
		b"0000000000000010000000",
		b"0000000000000001010010",
		b"0000000000000000100011",
		b"1111111111111111110101",
		b"1111111111111111000101",
		b"1111111111111110010110",
		b"1111111111111101100101",
		b"1111111111111100110101",
		b"1111111111111100000100",
		b"1111111111111011010011",
		b"1111111111111010100001",
		b"1111111111111001110000",
		b"1111111111111000111101",
		b"1111111111111000001011",
		b"1111111111110111011000",
		b"1111111111110110100110",
		b"1111111111110101110010",
		b"1111111111110100111111",
		b"1111111111110100001100",
		b"1111111111110011011000",
		b"1111111111110010100100",
		b"1111111111110001110001",
		b"1111111111110000111101",
		b"1111111111110000001001",
		b"1111111111101111010100",
		b"1111111111101110100000",
		b"1111111111101101101100",
		b"1111111111101100111000",
		b"1111111111101100000100",
		b"1111111111101011010000",
		b"1111111111101010011100",
		b"1111111111101001101000",
		b"1111111111101000110100",
		b"1111111111101000000000",
		b"1111111111100111001100",
		b"1111111111100110011001",
		b"1111111111100101100110",
		b"1111111111100100110010",
		b"1111111111100011111111",
		b"1111111111100011001101",
		b"1111111111100010011010",
		b"1111111111100001101000",
		b"1111111111100000110110",
		b"1111111111100000000100",
		b"1111111111011111010011",
		b"1111111111011110100010",
		b"1111111111011101110001",
		b"1111111111011101000001",
		b"1111111111011100010001",
		b"1111111111011011100001",
		b"1111111111011010110010",
		b"1111111111011010000011",
		b"1111111111011001010100",
		b"1111111111011000100110",
		b"1111111111010111111001",
		b"1111111111010111001100",
		b"1111111111010110011111",
		b"1111111111010101110011",
		b"1111111111010101001000",
		b"1111111111010100011101",
		b"1111111111010011110011",
		b"1111111111010011001001",
		b"1111111111010010011111",
		b"1111111111010001110111",
		b"1111111111010001001111",
		b"1111111111010000100111",
		b"1111111111010000000000",
		b"1111111111001111011010",
		b"1111111111001110110100",
		b"1111111111001110001111",
		b"1111111111001101101011",
		b"1111111111001101001000",
		b"1111111111001100100101",
		b"1111111111001100000010",
		b"1111111111001011100001",
		b"1111111111001011000000",
		b"1111111111001010100000",
		b"1111111111001010000001",
		b"1111111111001001100010",
		b"1111111111001001000100",
		b"1111111111001000100111",
		b"1111111111001000001011",
		b"1111111111000111101111",
		b"1111111111000111010100",
		b"1111111111000110111010",
		b"1111111111000110100001",
		b"1111111111000110001001",
		b"1111111111000101110001",
		b"1111111111000101011010",
		b"1111111111000101000100",
		b"1111111111000100101111",
		b"1111111111000100011011",
		b"1111111111000100000111",
		b"1111111111000011110100",
		b"1111111111000011100011",
		b"1111111111000011010010",
		b"1111111111000011000001",
		b"1111111111000010110010",
		b"1111111111000010100011",
		b"1111111111000010010110",
		b"1111111111000010001001",
		b"1111111111000001111101",
		b"1111111111000001110010",
		b"1111111111000001100111",
		b"1111111111000001011110",
		b"1111111111000001010101",
		b"1111111111000001001110",
		b"1111111111000001000111",
		b"1111111111000001000001",
		b"1111111111000000111011",
		b"1111111111000000110111",
		b"1111111111000000110100",
		b"1111111111000000110001",
		b"1111111111000000101111",
		b"1111111111000000101110",
		b"1111111111000000101110",
		b"1111111111000000101110",
		b"1111111111000000110000",
		b"1111111111000000110010",
		b"1111111111000000110101",
		b"1111111111000000111001",
		b"1111111111000000111110",
		b"1111111111000001000100",
		b"1111111111000001001010",
		b"1111111111000001010001",
		b"1111111111000001011001",
		b"1111111111000001100010",
		b"1111111111000001101011",
		b"1111111111000001110110",
		b"1111111111000010000001",
		b"1111111111000010001100",
		b"1111111111000010011001",
		b"1111111111000010100110",
		b"1111111111000010110100",
		b"1111111111000011000011",
		b"1111111111000011010011",
		b"1111111111000011100011",
		b"1111111111000011110100",
		b"1111111111000100000101",
		b"1111111111000100011000",
		b"1111111111000100101011",
		b"1111111111000100111110",
		b"1111111111000101010011",
		b"1111111111000101101000",
		b"1111111111000101111101",
		b"1111111111000110010011",
		b"1111111111000110101010",
		b"1111111111000111000010",
		b"1111111111000111011010",
		b"1111111111000111110011",
		b"1111111111001000001100",
		b"1111111111001000100110",
		b"1111111111001001000000",
		b"1111111111001001011011",
		b"1111111111001001110111",
		b"1111111111001010010011",
		b"1111111111001010110000",
		b"1111111111001011001101",
		b"1111111111001011101011",
		b"1111111111001100001001",
		b"1111111111001100100111",
		b"1111111111001101000110",
		b"1111111111001101100110",
		b"1111111111001110000110",
		b"1111111111001110100111",
		b"1111111111001111000111",
		b"1111111111001111101001",
		b"1111111111010000001010",
		b"1111111111010000101100",
		b"1111111111010001001111",
		b"1111111111010001110010",
		b"1111111111010010010101",
		b"1111111111010010111000",
		b"1111111111010011011100",
		b"1111111111010100000001",
		b"1111111111010100100101",
		b"1111111111010101001010",
		b"1111111111010101101111",
		b"1111111111010110010100",
		b"1111111111010110111010",
		b"1111111111010111100000",
		b"1111111111011000000110",
		b"1111111111011000101100",
		b"1111111111011001010011",
		b"1111111111011001111001",
		b"1111111111011010100000",
		b"1111111111011011000111",
		b"1111111111011011101111",
		b"1111111111011100010110",
		b"1111111111011100111110",
		b"1111111111011101100101",
		b"1111111111011110001101",
		b"1111111111011110110101",
		b"1111111111011111011101",
		b"1111111111100000000101",
		b"1111111111100000101110",
		b"1111111111100001010110",
		b"1111111111100001111110",
		b"1111111111100010100110",
		b"1111111111100011001111",
		b"1111111111100011110111",
		b"1111111111100100100000",
		b"1111111111100101001000",
		b"1111111111100101110001",
		b"1111111111100110011001",
		b"1111111111100111000001",
		b"1111111111100111101010",
		b"1111111111101000010010",
		b"1111111111101000111010",
		b"1111111111101001100010",
		b"1111111111101010001010",
		b"1111111111101010110010",
		b"1111111111101011011010",
		b"1111111111101100000010",
		b"1111111111101100101001",
		b"1111111111101101010001",
		b"1111111111101101111000",
		b"1111111111101110011111",
		b"1111111111101111000110",
		b"1111111111101111101101",
		b"1111111111110000010100",
		b"1111111111110000111011",
		b"1111111111110001100001",
		b"1111111111110010000111",
		b"1111111111110010101101",
		b"1111111111110011010011",
		b"1111111111110011111000",
		b"1111111111110100011101",
		b"1111111111110101000010",
		b"1111111111110101100111",
		b"1111111111110110001100",
		b"1111111111110110110000",
		b"1111111111110111010100",
		b"1111111111110111111000",
		b"1111111111111000011011",
		b"1111111111111000111110",
		b"1111111111111001100001",
		b"1111111111111010000100",
		b"1111111111111010100110",
		b"1111111111111011001000",
		b"1111111111111011101010",
		b"1111111111111100001011",
		b"1111111111111100101100",
		b"1111111111111101001100",
		b"1111111111111101101101",
		b"1111111111111110001101",
		b"1111111111111110101100",
		b"1111111111111111001100",
		b"1111111111111111101011",
		b"0000000000000000001001",
		b"0000000000000000100111",
		b"0000000000000001000101",
		b"0000000000000001100011",
		b"0000000000000010000000",
		b"0000000000000010011100",
		b"0000000000000010111001",
		b"0000000000000011010101",
		b"0000000000000011110000",
		b"0000000000000100001011",
		b"0000000000000100100110",
		b"0000000000000101000000",
		b"0000000000000101011010",
		b"0000000000000101110100",
		b"0000000000000110001101",
		b"0000000000000110100110",
		b"0000000000000110111110",
		b"0000000000000111010110",
		b"0000000000000111101110",
		b"0000000000001000000101",
		b"0000000000001000011100",
		b"0000000000001000110010",
		b"0000000000001001001000",
		b"0000000000001001011101",
		b"0000000000001001110010",
		b"0000000000001010000111",
		b"0000000000001010011011",
		b"0000000000001010101111",
		b"0000000000001011000010",
		b"0000000000001011010101",
		b"0000000000001011101000",
		b"0000000000001011111010",
		b"0000000000001100001100",
		b"0000000000001100011101",
		b"0000000000001100101110",
		b"0000000000001100111110",
		b"0000000000001101001111",
		b"0000000000001101011110",
		b"0000000000001101101101",
		b"0000000000001101111100",
		b"0000000000001110001011",
		b"0000000000001110011001",
		b"0000000000001110100110",
		b"0000000000001110110100",
		b"0000000000001111000000",
		b"0000000000001111001101",
		b"0000000000001111011001",
		b"0000000000001111100101",
		b"0000000000001111110000",
		b"0000000000001111111011",
		b"0000000000010000000101",
		b"0000000000010000001111",
		b"0000000000010000011001",
		b"0000000000010000100010",
		b"0000000000010000101011",
		b"0000000000010000110100",
		b"0000000000010000111100",
		b"0000000000010001000100",
		b"0000000000010001001011",
		b"0000000000010001010010",
		b"0000000000010001011001",
		b"0000000000010001011111",
		b"0000000000010001100101",
		b"0000000000010001101011",
		b"0000000000010001110000",
		b"0000000000010001110101",
		b"0000000000010001111010",
		b"0000000000010001111110",
		b"0000000000010010000010",
		b"0000000000010010000110",
		b"0000000000010010001001",
		b"0000000000010010001100",
		b"0000000000010010001111",
		b"0000000000010010010010",
		b"0000000000010010010100",
		b"0000000000010010010101",
		b"0000000000010010010111",
		b"0000000000010010011000",
		b"0000000000010010011001",
		b"0000000000010010011010",
		b"0000000000010010011010",
		b"0000000000010010011010",
		b"0000000000010010011010",
		b"0000000000010010011001",
		b"0000000000010010011001",
		b"0000000000010010011000",
		b"0000000000010010010110",
		b"0000000000010010010101",
		b"0000000000010010010011",
		b"0000000000010010010001",
		b"0000000000010010001111",
		b"0000000000010010001100",
		b"0000000000010010001001",
		b"0000000000010010000111",
		b"0000000000010010000011",
		b"0000000000010010000000",
		b"0000000000010001111100",
		b"0000000000010001111001",
		b"0000000000010001110101",
		b"0000000000010001110000",
		b"0000000000010001101100",
		b"0000000000010001100111",
		b"0000000000010001100011",
		b"0000000000010001011110",
		b"0000000000010001011000",
		b"0000000000010001010011",
		b"0000000000010001001110",
		b"0000000000010001001000",
		b"0000000000010001000010",
		b"0000000000010000111100",
		b"0000000000010000110110",
		b"0000000000010000110000",
		b"0000000000010000101010",
		b"0000000000010000100011",
		b"0000000000010000011100",
		b"0000000000010000010110",
		b"0000000000010000001111",
		b"0000000000010000001000",
		b"0000000000010000000000",
		b"0000000000001111111001",
		b"0000000000001111110010",
		b"0000000000001111101010",
		b"0000000000001111100011",
		b"0000000000001111011011",
		b"0000000000001111010011",
		b"0000000000001111001011",
		b"0000000000001111000011",
		b"0000000000001110111011",
		b"0000000000001110110011",
		b"0000000000001110101011",
		b"0000000000001110100011",
		b"0000000000001110011011",
		b"0000000000001110010010",
		b"0000000000001110001010",
		b"0000000000001110000001",
		b"0000000000001101111001",
		b"0000000000001101110000",
		b"0000000000001101101000",
		b"0000000000001101011111",
		b"0000000000001101010110",
		b"0000000000001101001101",
		b"0000000000001101000101",
		b"0000000000001100111100",
		b"0000000000001100110011",
		b"0000000000001100101010",
		b"0000000000001100100001",
		b"0000000000001100011000",
		b"0000000000001100010000",
		b"0000000000001100000111",
		b"0000000000001011111110",
		b"0000000000001011110101",
		b"0000000000001011101100",
		b"0000000000001011100011",
		b"0000000000001011011010",
		b"0000000000001011010001",
		b"0000000000001011001000",
		b"0000000000001010111111",
		b"0000000000001010110110",
		b"0000000000001010101110",
		b"0000000000001010100101",
		b"0000000000001010011100",
		b"0000000000001010010011",
		b"0000000000001010001010",
		b"0000000000001010000001",
		b"0000000000001001111001",
		b"0000000000001001110000",
		b"0000000000001001100111",
		b"0000000000001001011111",
		b"0000000000001001010110",
		b"0000000000001001001110",
		b"0000000000001001000101",
		b"0000000000001000111101",
		b"0000000000001000110100",
		b"0000000000001000101100",
		b"0000000000001000100100",
		b"0000000000001000011011",
		b"0000000000001000010011",
		b"0000000000001000001011",
		b"0000000000001000000011",
		b"0000000000000111111011",
		b"0000000000000111110011",
		b"0000000000000111101011",
		b"0000000000000111100011",
		b"0000000000000111011011",
		b"0000000000000111010011",
		b"0000000000000111001011",
		b"0000000000000111000100",
		b"0000000000000110111100",
		b"0000000000000110110101",
		b"0000000000000110101101",
		b"0000000000000110100110",
		b"0000000000000110011110",
		b"0000000000000110010111",
		b"0000000000000110010000",
		b"0000000000000110001001",
		b"0000000000000110000010",
		b"0000000000000101111011",
		b"0000000000000101110100",
		b"0000000000000101101101",
		b"0000000000000101100110",
		b"0000000000000101100000",
		b"0000000000000101011001",
		b"0000000000000101010010",
		b"0000000000000101001100",
		b"0000000000000101000110",
		b"0000000000000100111111",
		b"0000000000000100111001",
		b"0000000000000100110011",
		b"0000000000000100101101",
		b"0000000000000100100111",
		b"0000000000000100100001",
		b"0000000000000100011011",
		b"0000000000000100010101",
		b"0000000000000100001111",
		b"0000000000000100001010",
		b"0000000000000100000100",
		b"0000000000000011111111",
		b"0000000000000011111001",
		b"0000000000000011110100",
		b"0000000000000011101111",
		b"0000000000000011101010",
		b"0000000000000011100100",
		b"0000000000000011011111",
		b"0000000000000011011010",
		b"0000000000000011010110",
		b"0000000000000011010001",
		b"0000000000000011001100",
		b"0000000000000011000111",
		b"0000000000000011000011",
		b"0000000000000010111110",
		b"0000000000000010111010",
		b"0000000000000010110101",
		b"0000000000000010110001",
		b"0000000000000010101101",
		b"0000000000000010101001",
		b"0000000000000010100101",
		b"0000000000000010100001",
		b"0000000000000010011101",
		b"0000000000000010011001",
		b"0000000000000010010101",
		b"0000000000000010010001",
		b"0000000000000010001110",
		b"0000000000000010001010",
		b"0000000000000010000111",
		b"0000000000000010000011",
		b"0000000000000010000000",
		b"0000000000000001111100",
		b"0000000000000001111001",
		b"0000000000000001110110",
		b"0000000000000001110011",
		b"0000000000000001110000",
		b"0000000000000001101101",
		b"0000000000000001101010",
		b"0000000000000001100111",
		b"0000000000000001100100",
		b"0000000000000001100001",
		b"0000000000000001011110",
		b"0000000000000001011100",
		b"0000000000000001011001",
		b"0000000000000001010110",
		b"0000000000000001010100",
		b"0000000000000001010010",
		b"0000000000000001001111",
		b"0000000000000001001101",
		b"0000000000000001001010",
		b"0000000000000001001000",
		b"0000000000000001000110",
		b"0000000000000001000100",
		b"0000000000000001000010",
		b"0000000000000001000000",
		b"0000000000000000111110",
		b"0000000000000000111100",
		b"0000000000000000111010",
		b"0000000000000000111000",
		b"0000000000000000110110",
		b"0000000000000000110101",
		b"0000000000000000110011",
		b"0000000000000000110001",
		b"0000000000000000110000",
		b"0000000000000000101110",
		b"0000000000000000101100",
		b"0000000000000000101011",
		b"0000000000000000101001",
		b"0000000000000000101000",
		b"0000000000000000100111",
		b"0000000000000000100101",
		b"0000000000000000100100",
		b"0000000000000000100011",
		b"0000000000000000100001",
		b"0000000000000000100000",
		b"0000000000000000011111",
		b"0000000000000000011110",
		b"0000000000000000011101",
		b"0000000000000000011100",
		b"0000000000000000011011",
		b"0000000000000000011010",
		b"0000000000000000011001",
		b"0000000000000000011000",
		b"0000000000000000010111",
		b"0000000000000000010110",
		b"0000000000000000010101",
		b"0000000000000000010100",
		b"0000000000000000010011",
		b"0000000000000000010011",
		b"0000000000000000010010",
		b"0000000000000000010001",
		b"0000000000000000010000",
		b"0000000000000000010000",
		b"0000000000000000001111",
		b"0000000000000000001110",
		b"0000000000000000001110",
		b"0000000000000000001101",
		b"0000000000000000001101",
		b"0000000000000000001100",
		b"0000000000000000001011",
		b"0000000000000000001011",
		b"0000000000000000001010",
		b"0000000000000000001010",
		b"0000000000000000001001",
		b"0000000000000000001001",
		b"0000000000000000001001",
		b"0000000000000000001000",
		b"0000000000000000001000",
		b"0000000000000000000111",
		b"0000000000000000000111",
		b"0000000000000000000111",
		b"0000000000000000000110",
		b"0000000000000000000110",
		b"0000000000000000000110",
		b"0000000000000000000101",
		b"0000000000000000000101",
		b"0000000000000000000101",
		b"0000000000000000000101",
		b"0000000000000000000100",
		b"0000000000000000000100",
		b"0000000000000000000100",
		b"0000000000000000000100",
		b"0000000000000000000011",
		b"0000000000000000000011",
		b"0000000000000000000011",
		b"0000000000000000000011",
		b"0000000000000000000011",
		b"0000000000000000000010",
		b"0000000000000000000010",
		b"0000000000000000000010",
		b"0000000000000000000010",
		b"0000000000000000000010",
		b"0000000000000000000010",
		b"0000000000000000000010",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000001",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000",
		b"0000000000000000000000"
	);

end src_rom_pkg;