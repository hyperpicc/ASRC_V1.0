library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package src_rom_pkg is

	constant COE_WIDTH	: integer := 26;
	constant COE_CENTRE	: signed( 25 downto 0 ) := b"01111111010111000010100100";

	type COE_ROM_TYPE is array( 4095 downto 0 ) of signed( 25 downto 0 );
	constant COE_ROM	 : COE_ROM_TYPE := (
		b"01111111010110010001010110",
		b"01111111010011111101101101",
		b"01111111010000000111101011",
		b"01111111001010101111010111",
		b"01111111000011110100111000",
		b"01111110111011011000010111",
		b"01111110110001011010000001",
		b"01111110100101111010000011",
		b"01111110011000111000101101",
		b"01111110001010010110010001",
		b"01111101111010010011000101",
		b"01111101101000101111011101",
		b"01111101010101101011110011",
		b"01111101000001001000100001",
		b"01111100101011000110000100",
		b"01111100010011100100111010",
		b"01111011111010100101100100",
		b"01111011100000001000100101",
		b"01111011000100001110100010",
		b"01111010100110111000000010",
		b"01111010001000000101101100",
		b"01111001100111111000001101",
		b"01111001000110010000010001",
		b"01111000100011001110100110",
		b"01110111111110110011111110",
		b"01110111011001000001001010",
		b"01110110110001110110111111",
		b"01110110001001010110010011",
		b"01110101011111011111111110",
		b"01110100110100010100111011",
		b"01110100000111110110000100",
		b"01110011011010000100010111",
		b"01110010101011000000110101",
		b"01110001111010101100011100",
		b"01110001001001001000010000",
		b"01110000010110010101010110",
		b"01101111100010010100110010",
		b"01101110101101000111101101",
		b"01101101110110101111010000",
		b"01101100111111001100100101",
		b"01101100000110100000111000",
		b"01101011001100101101010111",
		b"01101010010001110011010001",
		b"01101001010101110011110111",
		b"01101000011000110000011011",
		b"01100111011010101010001111",
		b"01100110011011100010101000",
		b"01100101011011011010111101",
		b"01100100011010010100100100",
		b"01100011011000010000110110",
		b"01100010010101010001001100",
		b"01100001010001010111000001",
		b"01100000001100100011110001",
		b"01011111000110111000111001",
		b"01011110000000010111110110",
		b"01011100111001000010001000",
		b"01011011110000111001001110",
		b"01011010100111111110101010",
		b"01011001011110010011111100",
		b"01011000010011111010101001",
		b"01010111001000110100010010",
		b"01010101111101000010011101",
		b"01010100110000100110101101",
		b"01010011100011100010101010",
		b"01010010010101110111110111",
		b"01010001000111100111111111",
		b"01001111111000110100100110",
		b"01001110101001011111010101",
		b"01001101011001101001110101",
		b"01001100001001010101101110",
		b"01001010111000100100101010",
		b"01001001100111011000010011",
		b"01001000010101110010010010",
		b"01000111000011110100010001",
		b"01000101110001011111111100",
		b"01000100011110110110111101",
		b"01000011001011111010111110",
		b"01000001111000101101101100",
		b"01000000100101010000110000",
		b"00111111010001100101110110",
		b"00111101111101101110101001",
		b"00111100101001101100110101",
		b"00111011010101100010000011",
		b"00111010000001001111111111",
		b"00111000101100111000010100",
		b"00110111011000011100101011",
		b"00110110000011111110110000",
		b"00110100101111100000001011",
		b"00110011011011000010101000",
		b"00110010000110100111101101",
		b"00110000110010010001000110",
		b"00101111011110000000011001",
		b"00101110001001110111001111",
		b"00101100110101110111001110",
		b"00101011100010000001111110",
		b"00101010001110011001000101",
		b"00101000111010111110000111",
		b"00100111100111110010101011",
		b"00100110010100111000010011",
		b"00100101000010010000100011",
		b"00100011101111111100111110",
		b"00100010011101111111000101",
		b"00100001001100011000011001",
		b"00011111111011001010011001",
		b"00011110101010010110100101",
		b"00011101011001111110011011",
		b"00011100001010000011010111",
		b"00011010111010100110110110",
		b"00011001101011101010010010",
		b"00011000011101001111000100",
		b"00010111001111010110100110",
		b"00010110000010000010001110",
		b"00010100110101010011010100",
		b"00010011101001001011001011",
		b"00010010011101101011000111",
		b"00010001010010110100011100",
		b"00010000001000101000011001",
		b"00001110111111001000001110",
		b"00001101110110010101001011",
		b"00001100101110010000011011",
		b"00001011100110111011001011",
		b"00001010100000010110100011",
		b"00001001011010100011101110",
		b"00001000010101100011110001",
		b"00000111010001010111110010",
		b"00000110001110000000110110",
		b"00000101001011011111111110",
		b"00000100001001110110001100",
		b"00000011001001000100011101",
		b"00000010001001001011110010",
		b"00000001001010001101000101",
		b"00000000001100001001001111",
		b"11111111001111000001001010",
		b"11111110010010110101101101",
		b"11111101010111100111101100",
		b"11111100011101010111111011",
		b"11111011100100000111001100",
		b"11111010101011110110001110",
		b"11111001110100100101110000",
		b"11111000111110010110011101",
		b"11111000001001001001000000",
		b"11110111010100111110000011",
		b"11110110100001110110001011",
		b"11110101101111110001111110",
		b"11110100111110110001111110",
		b"11110100001110110110101110",
		b"11110011100000000000101100",
		b"11110010110010010000010111",
		b"11110010000101100110001001",
		b"11110001011010000010011110",
		b"11110000101111100101101100",
		b"11110000000110010000001010",
		b"11101111011110000010001101",
		b"11101110110110111100000110",
		b"11101110010000111110000110",
		b"11101101101100001000011100",
		b"11101101001000011011010101",
		b"11101100100101110110111011",
		b"11101100000100011011010111",
		b"11101011100100001000110010",
		b"11101011000100111111001110",
		b"11101010100110111110110010",
		b"11101010001010000111011110",
		b"11101001101110011001010001",
		b"11101001010011110100001010",
		b"11101000111010011000000101",
		b"11101000100010000100111011",
		b"11101000001010111010100111",
		b"11100111110100111000111101",
		b"11100111011111111111110100",
		b"11100111001100001110111110",
		b"11100110111001100110001101",
		b"11100110101000000101010000",
		b"11100110010111101011110110",
		b"11100110001000011001101010",
		b"11100101111010001110010111",
		b"11100101101101001001100110",
		b"11100101100001001010111110",
		b"11100101010110010010000100",
		b"11100101001100011110011101",
		b"11100101000011101111101010",
		b"11100100111100000101001101",
		b"11100100110101011110100100",
		b"11100100101111111011001110",
		b"11100100101011011010100110",
		b"11100100100111111100000110",
		b"11100100100101011111001001",
		b"11100100100100000011000101",
		b"11100100100011100111010000",
		b"11100100100100001011000000",
		b"11100100100101101101101000",
		b"11100100101000001110011010",
		b"11100100101011101100100101",
		b"11100100110000000111011100",
		b"11100100110101011110001011",
		b"11100100111011101111111110",
		b"11100101000010111100000011",
		b"11100101001011000001100010",
		b"11100101010011111111100110",
		b"11100101011101110101010110",
		b"11100101101000100001111010",
		b"11100101110100000100011000",
		b"11100110000000011011110101",
		b"11100110001101100111010100",
		b"11100110011011100101111000",
		b"11100110101010010110100100",
		b"11100110111001111000011001",
		b"11100111001010001010010110",
		b"11100111011011001011011011",
		b"11100111101100111010100111",
		b"11100111111111010110110111",
		b"11101000010010011111001000",
		b"11101000100110010010010110",
		b"11101000111010101111011101",
		b"11101001001111110101011000",
		b"11101001100101100011000001",
		b"11101001111011110111010001",
		b"11101010010010110001000010",
		b"11101010101010001111001101",
		b"11101011000010010000101000",
		b"11101011011010110100001101",
		b"11101011110011111000110001",
		b"11101100001101011101001100",
		b"11101100100111100000010101",
		b"11101101000010000001000000",
		b"11101101011100111110000110",
		b"11101101111000010110011010",
		b"11101110010100001000110011",
		b"11101110110000010100000100",
		b"11101111001100110111000100",
		b"11101111101001110000101000",
		b"11110000000110111111100011",
		b"11110000100100100010101100",
		b"11110001000010011000110110",
		b"11110001100000100000110111",
		b"11110001111110111001100100",
		b"11110010011101100001110001",
		b"11110010111100011000010100",
		b"11110011011011011100000001",
		b"11110011111010101011101111",
		b"11110100011010000110010010",
		b"11110100111001101010100001",
		b"11110101011001010111010010",
		b"11110101111001001011011011",
		b"11110110011001000101110100",
		b"11110110111001000101010011",
		b"11110111011001001000110000",
		b"11110111111001001111000011",
		b"11111000011001010111000101",
		b"11111000111001011111101111",
		b"11111001011001100111111010",
		b"11111001111001101110100001",
		b"11111010011001110010011101",
		b"11111010111001110010101100",
		b"11111011011001101110001000",
		b"11111011111001100011101110",
		b"11111100011001010010011011",
		b"11111100111000111001001111",
		b"11111101011000010111000110",
		b"11111101110111101011000010",
		b"11111110010110110100000010",
		b"11111110110101110001001000",
		b"11111111010100100001010110",
		b"11111111110011000011101111",
		b"00000000010001010111010110",
		b"00000000101111011011010001",
		b"00000001001101001110100110",
		b"00000001101010110000011010",
		b"00000010000111111111110110",
		b"00000010100100111100000010",
		b"00000011000001100100001000",
		b"00000011011101110111010011",
		b"00000011111001110100101111",
		b"00000100010101011011101001",
		b"00000100110000101011001110",
		b"00000101001011100010101111",
		b"00000101100110000001011010",
		b"00000110000000000110100010",
		b"00000110011001110001011001",
		b"00000110110011000001010011",
		b"00000111001011110101100110",
		b"00000111100100001101100110",
		b"00000111111100001000101100",
		b"00001000010011100110010000",
		b"00001000101010100101101101",
		b"00001001000001000110011100",
		b"00001001010111000111111100",
		b"00001001101100101001101001",
		b"00001010000001101011000010",
		b"00001010010110001011101000",
		b"00001010101010001010111101",
		b"00001010111101101000100010",
		b"00001011010000100011111101",
		b"00001011100010111100110011",
		b"00001011110100110010101011",
		b"00001100000110000101001100",
		b"00001100010110110100000001",
		b"00001100100110111110110100",
		b"00001100110110100101010010",
		b"00001101000101100111001000",
		b"00001101010100000100000100",
		b"00001101100001111011111000",
		b"00001101101111001110010100",
		b"00001101111011111011001011",
		b"00001110001000000010010011",
		b"00001110010011100011011111",
		b"00001110011110011110101000",
		b"00001110101000110011100101",
		b"00001110110010100010010001",
		b"00001110111011101010100101",
		b"00001111000100001100011110",
		b"00001111001100000111111001",
		b"00001111010011011100110110",
		b"00001111011010001011010100",
		b"00001111100000010011010101",
		b"00001111100101110100111011",
		b"00001111101010110000001011",
		b"00001111101111000101001010",
		b"00001111110010110011111101",
		b"00001111110101111100101101",
		b"00001111111000011111100100",
		b"00001111111010011100101001",
		b"00001111111011110100001010",
		b"00001111111100100110010011",
		b"00001111111100110011010001",
		b"00001111111100011011010100",
		b"00001111111011011110101011",
		b"00001111111001111101101000",
		b"00001111110111111000011100",
		b"00001111110101001111011100",
		b"00001111110010000010111100",
		b"00001111101110010011010001",
		b"00001111101010000000110010",
		b"00001111100101001011110111",
		b"00001111011111110100111000",
		b"00001111011001111100001111",
		b"00001111010011100010010111",
		b"00001111001100100111101100",
		b"00001111000101001100101010",
		b"00001110111101010001101110",
		b"00001110110100110111010111",
		b"00001110101011111110000101",
		b"00001110100010100110010110",
		b"00001110011000110000101110",
		b"00001110001110011101101100",
		b"00001110000011101101110101",
		b"00001101111000100001101011",
		b"00001101101100111001110010",
		b"00001101100000110110110000",
		b"00001101010100011001001010",
		b"00001101000111100001100110",
		b"00001100111010010000101010",
		b"00001100101100100111000001",
		b"00001100011110100101001111",
		b"00001100010000001100000000",
		b"00001100000001011011111011",
		b"00001011110010010101101100",
		b"00001011100010111001111011",
		b"00001011010011001001010101",
		b"00001011000011000100100101",
		b"00001010110010101100010110",
		b"00001010100010000001010100",
		b"00001010010001000100001101",
		b"00001001111111110101101101",
		b"00001001101110010110100001",
		b"00001001011100100111010111",
		b"00001001001010101000111110",
		b"00001000111000011100000010",
		b"00001000100110000001010011",
		b"00001000010011011001011111",
		b"00001000000000100101010101",
		b"00000111101101100101100100",
		b"00000111011010011010111011",
		b"00000111000111000110001001",
		b"00000110110011100111111110",
		b"00000110100000000001001000",
		b"00000110001100010010011000",
		b"00000101111000011100011101",
		b"00000101100100100000000101",
		b"00000101010000011110000010",
		b"00000100111100010111000000",
		b"00000100101000001011110001",
		b"00000100010011111101000011",
		b"00000011111111101011100100",
		b"00000011101011011000000101",
		b"00000011010111000011010010",
		b"00000011000010101101111100",
		b"00000010101110011000101111",
		b"00000010011010000100011010",
		b"00000010000101110001101010",
		b"00000001110001100001001110",
		b"00000001011101010011110001",
		b"00000001001001001010000000",
		b"00000000110101000100101000",
		b"00000000100001000100010101",
		b"00000000001101001001110010",
		b"11111111111001010101101010",
		b"11111111100101101000100111",
		b"11111111010010000011010101",
		b"11111110111110100110011101",
		b"11111110101011010010100111",
		b"11111110011000001000011100",
		b"11111110000101001000100101",
		b"11111101110010010011101001",
		b"11111101011111101010001111",
		b"11111101001101001100111101",
		b"11111100111010111100011001",
		b"11111100101000111001001000",
		b"11111100010111000011101110",
		b"11111100000101011100101111",
		b"11111011110100000100101110",
		b"11111011100010111100001110",
		b"11111011010010000011110000",
		b"11111011000001011011110101",
		b"11111010110001000100111101",
		b"11111010100000111111101000",
		b"11111010010001001100010100",
		b"11111010000001101011100000",
		b"11111001110010011101100111",
		b"11111001100011100011000111",
		b"11111001010100111100011011",
		b"11111001000110101001111101",
		b"11111000111000101100000111",
		b"11111000101011000011010011",
		b"11111000011101101111111000",
		b"11111000010000110010001110",
		b"11111000000100001010101010",
		b"11110111110111111001100010",
		b"11110111101011111111001100",
		b"11110111100000011011111010",
		b"11110111010101001111111111",
		b"11110111001010011011101101",
		b"11110110111111111111010110",
		b"11110110110101111011001001",
		b"11110110101100001111010100",
		b"11110110100010111100001000",
		b"11110110011010000001110000",
		b"11110110010001100000011001",
		b"11110110001001011000001110",
		b"11110110000001101001011010",
		b"11110101111010010100000111",
		b"11110101110011011000011101",
		b"11110101101100110110100011",
		b"11110101100110101110100001",
		b"11110101100001000000011100",
		b"11110101011011101100011000",
		b"11110101010110110010011011",
		b"11110101010010010010100111",
		b"11110101001110001100111101",
		b"11110101001010100001100000",
		b"11110101000111010000001111",
		b"11110101000100011001001001",
		b"11110101000001111100001110",
		b"11110100111111111001011010",
		b"11110100111110010000101010",
		b"11110100111101000001111001",
		b"11110100111100001101000011",
		b"11110100111011110010000010",
		b"11110100111011110000101101",
		b"11110100111100001000111111",
		b"11110100111100111010101101",
		b"11110100111110000101101111",
		b"11110100111111101001111010",
		b"11110101000001100111000010",
		b"11110101000011111100111100",
		b"11110101000110101011011011",
		b"11110101001001110010010001",
		b"11110101001101010001010000",
		b"11110101010001001000001001",
		b"11110101010101010110101011",
		b"11110101011001111100100101",
		b"11110101011110111001101000",
		b"11110101100100001101011111",
		b"11110101101001110111111000",
		b"11110101101111111000100000",
		b"11110101110110001111000011",
		b"11110101111100111011001010",
		b"11110110000011111100100001",
		b"11110110001011010010110001",
		b"11110110010010111101100100",
		b"11110110011010111100100001",
		b"11110110100011001111010001",
		b"11110110101011110101011011",
		b"11110110110100101110100101",
		b"11110110111101111010010110",
		b"11110111000111011000010011",
		b"11110111010001001000000010",
		b"11110111011011001001000110",
		b"11110111100101011011000101",
		b"11110111101111111101100001",
		b"11110111111010101111111110",
		b"11111000000101110001111111",
		b"11111000010001000011000101",
		b"11111000011100100010110011",
		b"11111000101000010000101011",
		b"11111000110100001100001101",
		b"11111001000000010100111010",
		b"11111001001100101010010011",
		b"11111001011001001011111001",
		b"11111001100101111001001010",
		b"11111001110010110001100111",
		b"11111001111111110100101110",
		b"11111010001101000010000001",
		b"11111010011010011000111100",
		b"11111010100111111000111111",
		b"11111010110101100001101000",
		b"11111011000011010010010111",
		b"11111011010001001010101000",
		b"11111011011111001001111011",
		b"11111011101101001111101101",
		b"11111011111011011011011101",
		b"11111100001001101100101000",
		b"11111100011000000010101100",
		b"11111100100110011101000111",
		b"11111100110100111011011000",
		b"11111101000011011100111010",
		b"11111101010010000001001110",
		b"11111101100000100111110000",
		b"11111101101111001111111111",
		b"11111101111101111001011000",
		b"11111110001100100011011011",
		b"11111110011011001101100100",
		b"11111110101001110111010100",
		b"11111110111000100000000111",
		b"11111111000111000111011110",
		b"11111111010101101100110111",
		b"11111111100100001111110001",
		b"11111111110010101111101100",
		b"00000000000001001100000111",
		b"00000000001111100100100011",
		b"00000000011101111000011111",
		b"00000000101100000111011101",
		b"00000000111010010000111100",
		b"00000001001000010100011110",
		b"00000001010110010001100101",
		b"00000001100100000111110010",
		b"00000001110001110110101000",
		b"00000001111111011101101000",
		b"00000010001100111100010111",
		b"00000010011010010010010111",
		b"00000010100111011111001101",
		b"00000010110100100010011100",
		b"00000011000001011011101010",
		b"00000011001110001010011011",
		b"00000011011010101110010101",
		b"00000011100111000110111111",
		b"00000011110011010011111111",
		b"00000011111111010100111011",
		b"00000100001011001001011101",
		b"00000100010110110001001100",
		b"00000100100010001011110001",
		b"00000100101101011000110110",
		b"00000100111000011000000100",
		b"00000101000011001001000101",
		b"00000101001101101011100110",
		b"00000101010111111111010001",
		b"00000101100010000011110011",
		b"00000101101011111000111001",
		b"00000101110101011110010001",
		b"00000101111110110011101001",
		b"00000110000111111000101110",
		b"00000110010000101101010010",
		b"00000110011001010001000100",
		b"00000110100001100011110101",
		b"00000110101001100101010111",
		b"00000110110001010101011010",
		b"00000110111000110011110011",
		b"00000111000000000000010101",
		b"00000111000110111010110100",
		b"00000111001101100011000101",
		b"00000111010011111000111101",
		b"00000111011001111100010010",
		b"00000111011111101100111100",
		b"00000111100101001010110010",
		b"00000111101010010101101101",
		b"00000111101111001101100100",
		b"00000111110011110010010100",
		b"00000111111000000011110100",
		b"00000111111100000010000010",
		b"00000111111111101100111000",
		b"00001000000011000100010100",
		b"00001000000110001000010001",
		b"00001000001000111000110000",
		b"00001000001011010101101101",
		b"00001000001101011111001000",
		b"00001000001111010101000010",
		b"00001000010000110111011100",
		b"00001000010010000110010101",
		b"00001000010011000001110010",
		b"00001000010011101001110100",
		b"00001000010011111110011111",
		b"00001000010011111111110111",
		b"00001000010011101110000001",
		b"00001000010011001001000010",
		b"00001000010010010001000001",
		b"00001000010001000110000100",
		b"00001000001111101000010100",
		b"00001000001101110111110111",
		b"00001000001011110100110110",
		b"00001000001001011111011011",
		b"00001000000110110111110001",
		b"00001000000011111110000000",
		b"00001000000000110010010110",
		b"00000111111101010100111100",
		b"00000111111001100110000000",
		b"00000111110101100101101111",
		b"00000111110001010100010110",
		b"00000111101100110010000011",
		b"00000111100111111111000101",
		b"00000111100010111011101010",
		b"00000111011101101000000011",
		b"00000111011000000100100000",
		b"00000111010010010001010001",
		b"00000111001100001110100111",
		b"00000111000101111100110101",
		b"00000110111111011100001011",
		b"00000110111000101100111110",
		b"00000110110001101111011111",
		b"00000110101010100100000011",
		b"00000110100011001010111101",
		b"00000110011011100100100001",
		b"00000110010011110001000100",
		b"00000110001011110000111100",
		b"00000110000011100100011101",
		b"00000101111011001011111110",
		b"00000101110010100111110100",
		b"00000101101001111000010111",
		b"00000101100000111101111100",
		b"00000101010111111000111011",
		b"00000101001110101001101100",
		b"00000101000101010000100110",
		b"00000100111011101110000001",
		b"00000100110010000010010101",
		b"00000100101000001101111010",
		b"00000100011110010001001010",
		b"00000100010100001100011101",
		b"00000100001010000000001100",
		b"00000011111111101100110000",
		b"00000011110101010010100011",
		b"00000011101010110001111110",
		b"00000011100000001011011011",
		b"00000011010101011111010011",
		b"00000011001010101110000001",
		b"00000010111111110111111110",
		b"00000010110100111101100101",
		b"00000010101001111111001111",
		b"00000010011110111101010111",
		b"00000010010011111000010110",
		b"00000010001000110000101000",
		b"00000001111101100110100101",
		b"00000001110010011010101001",
		b"00000001100111001101001110",
		b"00000001011011111110101101",
		b"00000001010000101111100000",
		b"00000001000101100000000010",
		b"00000000111010010000101101",
		b"00000000101111000001111001",
		b"00000000100011110100000010",
		b"00000000011000100111011111",
		b"00000000001101011100101100",
		b"00000000000010010100000000",
		b"11111111110111001101110110",
		b"11111111101100001010100110",
		b"11111111100001001010101000",
		b"11111111010110001110010110",
		b"11111111001011010110000110",
		b"11111111000000100010010011",
		b"11111110110101110011010011",
		b"11111110101011001001011101",
		b"11111110100000100101001010",
		b"11111110010110000110101111",
		b"11111110001011101110100101",
		b"11111110000001011101000001",
		b"11111101110111010010011000",
		b"11111101101101001111000010",
		b"11111101100011010011010100",
		b"11111101011001011111100001",
		b"11111101001111110100000000",
		b"11111101000110010001000101",
		b"11111100111100110111000011",
		b"11111100110011100110001110",
		b"11111100101010011110111001",
		b"11111100100001100001010111",
		b"11111100011000101101111010",
		b"11111100010000000100110101",
		b"11111100000111100110011001",
		b"11111011111111010010110110",
		b"11111011110111001010011101",
		b"11111011101111001101011111",
		b"11111011100111011100001011",
		b"11111011011111110110110001",
		b"11111011011000011101011110",
		b"11111011010001010000100010",
		b"11111011001010010000001010",
		b"11111011000011011100100011",
		b"11111010111100110101111011",
		b"11111010110110011100011100",
		b"11111010110000010000010100",
		b"11111010101010010001101101",
		b"11111010100100100000110010",
		b"11111010011110111101101101",
		b"11111010011001101000100111",
		b"11111010010100100001101011",
		b"11111010001111101001000000",
		b"11111010001010111110101110",
		b"11111010000110100010111101",
		b"11111010000010010101110100",
		b"11111001111110010111011001",
		b"11111001111010100111110010",
		b"11111001110111000111000101",
		b"11111001110011110101010101",
		b"11111001110000110010101000",
		b"11111001101101111111000001",
		b"11111001101011011010100010",
		b"11111001101001000101010000",
		b"11111001100110111111001010",
		b"11111001100101001000010100",
		b"11111001100011100000101101",
		b"11111001100010001000010111",
		b"11111001100000111111010000",
		b"11111001100000000101011001",
		b"11111001011111011010110000",
		b"11111001011110111111010010",
		b"11111001011110110010111110",
		b"11111001011110110101110001",
		b"11111001011111000111101000",
		b"11111001011111101000011101",
		b"11111001100000011000001110",
		b"11111001100001010110110100",
		b"11111001100010100100001011",
		b"11111001100100000000001100",
		b"11111001100101101010110001",
		b"11111001100111100011110011",
		b"11111001101001101011001010",
		b"11111001101100000000101110",
		b"11111001101110100100010111",
		b"11111001110001010101111100",
		b"11111001110100010101010011",
		b"11111001110111100010010011",
		b"11111001111010111100110000",
		b"11111001111110100100100001",
		b"11111010000010011001011011",
		b"11111010000110011011010000",
		b"11111010001010101001110111",
		b"11111010001111000101000001",
		b"11111010010011101100100010",
		b"11111010011000100000001100",
		b"11111010011101011111110011",
		b"11111010100010101011000111",
		b"11111010101000000001111011",
		b"11111010101101100100000000",
		b"11111010110011010001000110",
		b"11111010111001001000111110",
		b"11111010111111001011011001",
		b"11111011000101011000000101",
		b"11111011001011101110110011",
		b"11111011010010001111010001",
		b"11111011011000111001010000",
		b"11111011011111101100011100",
		b"11111011100110101000100101",
		b"11111011101101101101011001",
		b"11111011110100111010100110",
		b"11111011111100001111111001",
		b"11111100000011101101000000",
		b"11111100001011010001100111",
		b"11111100010010111101011101",
		b"11111100011010110000001101",
		b"11111100100010101001100100",
		b"11111100101010101001001110",
		b"11111100110010101110111001",
		b"11111100111010111010010000",
		b"11111101000011001010111111",
		b"11111101001011100000110001",
		b"11111101010011111011010011",
		b"11111101011100011010010000",
		b"11111101100100111101010100",
		b"11111101101101100100001010",
		b"11111101110110001110011110",
		b"11111101111110111011111011",
		b"11111110000111101100001100",
		b"11111110010000011110111100",
		b"11111110011001010011110111",
		b"11111110100010001010101000",
		b"11111110101011000010111010",
		b"11111110110011111100011001",
		b"11111110111100110110101111",
		b"11111111000101110001101001",
		b"11111111001110101100110001",
		b"11111111010111100111110010",
		b"11111111100000100010011001",
		b"11111111101001011100010001",
		b"11111111110010010101000101",
		b"11111111111011001100100010",
		b"00000000000100000010010010",
		b"00000000001100110110000011",
		b"00000000010101100111100001",
		b"00000000011110010110010111",
		b"00000000100111000010010010",
		b"00000000101111101010111110",
		b"00000000111000010000001010",
		b"00000001000000110001100000",
		b"00000001001001001110110000",
		b"00000001010001100111100101",
		b"00000001011001111011101111",
		b"00000001100010001010111001",
		b"00000001101010010100110100",
		b"00000001110010011001001100",
		b"00000001111010010111110001",
		b"00000010000010010000010010",
		b"00000010001010000010011100",
		b"00000010010001101110000001",
		b"00000010011001010010101111",
		b"00000010100000110000010111",
		b"00000010101000000110101001",
		b"00000010101111010101010101",
		b"00000010110110011100001101",
		b"00000010111101011011000001",
		b"00000011000100010001100100",
		b"00000011001010111111100111",
		b"00000011010001100100111100",
		b"00000011011000000001010111",
		b"00000011011110010100101010",
		b"00000011100100011110101000",
		b"00000011101010011111000101",
		b"00000011110000010101110110",
		b"00000011110110000010101111",
		b"00000011111011100101100101",
		b"00000100000000111110001101",
		b"00000100000110001100011101",
		b"00000100001011010000001010",
		b"00000100010000001001001101",
		b"00000100010100110111011010",
		b"00000100011001011010101010",
		b"00000100011101110010110101",
		b"00000100100001111111110011",
		b"00000100100110000001011100",
		b"00000100101001110111101001",
		b"00000100101101100010010100",
		b"00000100110001000001010111",
		b"00000100110100010100101100",
		b"00000100110111011100001110",
		b"00000100111010010111111000",
		b"00000100111101000111100110",
		b"00000100111111101011010100",
		b"00000101000010000010111110",
		b"00000101000100001110100010",
		b"00000101000110001101111101",
		b"00000101001000000001001100",
		b"00000101001001101000001111",
		b"00000101001011000011000011",
		b"00000101001100010001101001",
		b"00000101001101010011111111",
		b"00000101001110001010000110",
		b"00000101001110110011111111",
		b"00000101001111010001101010",
		b"00000101001111100011001000",
		b"00000101001111101000011100",
		b"00000101001111100001101000",
		b"00000101001111001110101111",
		b"00000101001110101111110011",
		b"00000101001110000100111001",
		b"00000101001101001110000011",
		b"00000101001100001011010111",
		b"00000101001010111100111010",
		b"00000101001001100010110000",
		b"00000101000111111100111111",
		b"00000101000110001011101101",
		b"00000101000100001111000001",
		b"00000101000010000111000001",
		b"00000100111111110011110100",
		b"00000100111101010101100010",
		b"00000100111010101100010100",
		b"00000100110111111000010000",
		b"00000100110100111001100000",
		b"00000100110001110000001101",
		b"00000100101110011100100000",
		b"00000100101010111110100011",
		b"00000100100111010110100000",
		b"00000100100011100100100010",
		b"00000100011111101000110010",
		b"00000100011011100011011100",
		b"00000100010111010100101011",
		b"00000100010010111100101100",
		b"00000100001110011011101001",
		b"00000100001001110001101111",
		b"00000100000100111111001010",
		b"00000100000000000100001000",
		b"00000011111011000000110101",
		b"00000011110101110101011111",
		b"00000011110000100010010011",
		b"00000011101011000111011110",
		b"00000011100101100101010000",
		b"00000011011111111011110101",
		b"00000011011010001011011101",
		b"00000011010100010100010110",
		b"00000011001110010110101111",
		b"00000011001000010010110111",
		b"00000011000010001000111101",
		b"00000010111011111001010001",
		b"00000010110101100100000001",
		b"00000010101111001001011110",
		b"00000010101000101001111000",
		b"00000010100010000101011110",
		b"00000010011011011100100001",
		b"00000010010100101111010001",
		b"00000010001101111101111101",
		b"00000010000111001000110111",
		b"00000010000000010000001111",
		b"00000001111001010100010110",
		b"00000001110010010101011011",
		b"00000001101011010011110000",
		b"00000001100100001111100110",
		b"00000001011101001001001101",
		b"00000001010110000000110110",
		b"00000001001110110110110010",
		b"00000001000111101011010001",
		b"00000001000000011110100101",
		b"00000000111001010000111110",
		b"00000000110010000010101101",
		b"00000000101010110100000011",
		b"00000000100011100101010000",
		b"00000000011100010110100110",
		b"00000000010101001000010101",
		b"00000000001101111010101101",
		b"00000000000110101101111110",
		b"11111111111111100010011011",
		b"11111111111000011000010001",
		b"11111111110001001111110011",
		b"11111111101010001001001111",
		b"11111111100011000100110111",
		b"11111111011100000010111001",
		b"11111111010101000011100101",
		b"11111111001110000111001100",
		b"11111111000111001101111100",
		b"11111111000000011000000101",
		b"11111110111001100101110110",
		b"11111110110010110111011101",
		b"11111110101100001101001010",
		b"11111110100101100111001011",
		b"11111110011111000101101111",
		b"11111110011000101001000011",
		b"11111110010010010001010101",
		b"11111110001011111110110100",
		b"11111110000101110001101100",
		b"11111101111111101010001011",
		b"11111101111001101000011110",
		b"11111101110011101100110010",
		b"11111101101101110111010010",
		b"11111101101000001000001101",
		b"11111101100010011111101100",
		b"11111101011100111101111101",
		b"11111101010111100011001010",
		b"11111101010010001111011111",
		b"11111101001101000011000110",
		b"11111101000111111110001010",
		b"11111101000011000000110110",
		b"11111100111110001011010011",
		b"11111100111001011101101010",
		b"11111100110100111000000110",
		b"11111100110000011010101111",
		b"11111100101100000101101110",
		b"11111100100111111001001100",
		b"11111100100011110101001111",
		b"11111100011111111010000001",
		b"11111100011100000111101000",
		b"11111100011000011110001011",
		b"11111100010100111101110001",
		b"11111100010001100110100001",
		b"11111100001110011000100001",
		b"11111100001011010011110101",
		b"11111100001000011000100100",
		b"11111100000101100110110001",
		b"11111100000010111110100011",
		b"11111100000000011111111101",
		b"11111011111110001011000011",
		b"11111011111011111111111000",
		b"11111011111001111110100000",
		b"11111011111000000110111101",
		b"11111011110110011001010010",
		b"11111011110100110101100001",
		b"11111011110011011011101011",
		b"11111011110010001011110010",
		b"11111011110001000101110111",
		b"11111011110000001001111011",
		b"11111011101111010111111101",
		b"11111011101110101111111110",
		b"11111011101110010001111101",
		b"11111011101101111101111001",
		b"11111011101101110011110010",
		b"11111011101101110011100101",
		b"11111011101101111101010001",
		b"11111011101110010000110011",
		b"11111011101110101110001001",
		b"11111011101111010101010001",
		b"11111011110000000110000110",
		b"11111011110001000000100101",
		b"11111011110010000100101010",
		b"11111011110011010010010010",
		b"11111011110100101001010110",
		b"11111011110110001001110011",
		b"11111011110111110011100011",
		b"11111011111001100110100001",
		b"11111011111011100010100111",
		b"11111011111101100111101101",
		b"11111011111111110101101111",
		b"11111100000010001100100101",
		b"11111100000100101100001001",
		b"11111100000111010100010001",
		b"11111100001010000100111000",
		b"11111100001100111101110101",
		b"11111100001111111111000000",
		b"11111100010011001000010000",
		b"11111100010110011001011101",
		b"11111100011001110010011101",
		b"11111100011101010011000111",
		b"11111100100000111011010010",
		b"11111100100100101010110100",
		b"11111100101000100001100011",
		b"11111100101100011111010100",
		b"11111100110000100011111110",
		b"11111100110100101111010101",
		b"11111100111001000001001111",
		b"11111100111101011001100001",
		b"11111101000001110111111111",
		b"11111101000110011100011101",
		b"11111101001011000110110001",
		b"11111101001111110110101110",
		b"11111101010100101100001000",
		b"11111101011001100110110011",
		b"11111101011110100110100100",
		b"11111101100011101011001100",
		b"11111101101000110100100000",
		b"11111101101110000010010100",
		b"11111101110011010100011001",
		b"11111101111000101010100100",
		b"11111101111110000100100111",
		b"11111110000011100010010101",
		b"11111110001001000011100000",
		b"11111110001110100111111100",
		b"11111110010100001111011010",
		b"11111110011001111001101110",
		b"11111110011111100110101010",
		b"11111110100101010110000000",
		b"11111110101011000111100010",
		b"11111110110000111011000011",
		b"11111110110110110000010110",
		b"11111110111100100111001011",
		b"11111111000010011111010110",
		b"11111111001000011000101001",
		b"11111111001110010010110101",
		b"11111111010100001101101110",
		b"11111111011010001001000101",
		b"11111111100000000100101100",
		b"11111111100110000000010111",
		b"11111111101011111011110111",
		b"11111111110001110110111110",
		b"11111111110111110001100000",
		b"11111111111101101011001110",
		b"00000000000011100011111011",
		b"00000000001001011011011010",
		b"00000000001111010001011101",
		b"00000000010101000101110111",
		b"00000000011010111000011100",
		b"00000000100000101000111110",
		b"00000000100110010111010000",
		b"00000000101100000011000101",
		b"00000000110001101100010010",
		b"00000000110111010010101001",
		b"00000000111100110101111101",
		b"00000001000010010110000100",
		b"00000001000111110010110000",
		b"00000001001101001011110110",
		b"00000001010010100001001010",
		b"00000001010111110010100001",
		b"00000001011100111111101110",
		b"00000001100010001000101000",
		b"00000001100111001101000010",
		b"00000001101100001100110010",
		b"00000001110001000111101101",
		b"00000001110101111101101010",
		b"00000001111010101110011101",
		b"00000001111111011001111100",
		b"00000010000011111111111111",
		b"00000010001000100000011010",
		b"00000010001100111011000110",
		b"00000010010001001111111000",
		b"00000010010101011110101000",
		b"00000010011001100111001110",
		b"00000010011101101001100001",
		b"00000010100001100101011000",
		b"00000010100101011010101100",
		b"00000010101001001001010110",
		b"00000010101100110001001110",
		b"00000010110000010010001100",
		b"00000010110011101100001011",
		b"00000010110110111111000011",
		b"00000010111010001010101110",
		b"00000010111101001111000111",
		b"00000011000000001100000111",
		b"00000011000011000001101001",
		b"00000011000101101111101000",
		b"00000011001000010101111111",
		b"00000011001010110100101001",
		b"00000011001101001011100011",
		b"00000011001111011010101000",
		b"00000011010001100001110100",
		b"00000011010011100001000101",
		b"00000011010101011000010110",
		b"00000011010111000111100110",
		b"00000011011000101110110001",
		b"00000011011010001101110101",
		b"00000011011011100100110010",
		b"00000011011100110011100011",
		b"00000011011101111010001010",
		b"00000011011110111000100100",
		b"00000011011111101110110000",
		b"00000011100000011100101111",
		b"00000011100001000010100000",
		b"00000011100001100000000011",
		b"00000011100001110101011001",
		b"00000011100010000010100011",
		b"00000011100010000111100001",
		b"00000011100010000100010101",
		b"00000011100001111001000000",
		b"00000011100001100101100101",
		b"00000011100001001010000101",
		b"00000011100000100110100100",
		b"00000011011111111011000011",
		b"00000011011111000111100110",
		b"00000011011110001100010000",
		b"00000011011101001001000100",
		b"00000011011011111110001000",
		b"00000011011010101011011110",
		b"00000011011001010001001011",
		b"00000011010111101111010100",
		b"00000011010110000101111101",
		b"00000011010100010101001100",
		b"00000011010010011101000111",
		b"00000011010000011101110010",
		b"00000011001110010111010100",
		b"00000011001100001001110011",
		b"00000011001001110101010101",
		b"00000011000111011010000010",
		b"00000011000100110111111111",
		b"00000011000010001111010100",
		b"00000010111111100000001000",
		b"00000010111100101010100010",
		b"00000010111001101110101011",
		b"00000010110110101100101010",
		b"00000010110011100100101000",
		b"00000010110000010110101100",
		b"00000010101101000010111111",
		b"00000010101001101001101010",
		b"00000010100110001010110110",
		b"00000010100010100110101100",
		b"00000010011110111101010100",
		b"00000010011011001110111000",
		b"00000010010111011011100010",
		b"00000010010011100011011100",
		b"00000010001111100110101110",
		b"00000010001011100101100100",
		b"00000010000111100000000111",
		b"00000010000011010110100001",
		b"00000001111111001000111101",
		b"00000001111010110111100101",
		b"00000001110110100010100100",
		b"00000001110010001010000011",
		b"00000001101101101110001111",
		b"00000001101001001111010010",
		b"00000001100100101101010110",
		b"00000001100000001000100111",
		b"00000001011011100001001111",
		b"00000001010110110111011011",
		b"00000001010010001011010100",
		b"00000001001101011101000110",
		b"00000001001000101100111101",
		b"00000001000011111011000100",
		b"00000000111111000111100110",
		b"00000000111010010010101110",
		b"00000000110101011100101000",
		b"00000000110000100101011111",
		b"00000000101011101101011110",
		b"00000000100110110100110010",
		b"00000000100001111011100100",
		b"00000000011101000010000010",
		b"00000000011000001000010101",
		b"00000000010011001110101010",
		b"00000000001110010101001011",
		b"00000000001001011100000100",
		b"00000000000100100011100000",
		b"11111111111111101011101010",
		b"11111111111010110100101110",
		b"11111111110101111110110110",
		b"11111111110001001010001101",
		b"11111111101100010110111110",
		b"11111111100111100101010100",
		b"11111111100010110101011001",
		b"11111111011110000111011001",
		b"11111111011001011011011110",
		b"11111111010100110001110010",
		b"11111111010000001010011111",
		b"11111111001011100101110000",
		b"11111111000111000011101110",
		b"11111111000010100100100101",
		b"11111110111110001000011100",
		b"11111110111001101111011111",
		b"11111110110101011001110111",
		b"11111110110001000111101100",
		b"11111110101100111001001001",
		b"11111110101000101110010110",
		b"11111110100100100111011100",
		b"11111110100000100100100101",
		b"11111110011100100101111000",
		b"11111110011000101011011110",
		b"11111110010100110101011111",
		b"11111110010001000100000100",
		b"11111110001101010111010100",
		b"11111110001001101111010110",
		b"11111110000110001100010011",
		b"11111110000010101110010001",
		b"11111101111111010101011000",
		b"11111101111100000001101111",
		b"11111101111000110011011011",
		b"11111101110101101010100101",
		b"11111101110010100111010001",
		b"11111101101111101001100110",
		b"11111101101100110001101001",
		b"11111101101001111111100001",
		b"11111101100111010011010011",
		b"11111101100100101101000011",
		b"11111101100010001100110111",
		b"11111101011111110010110100",
		b"11111101011101011110111100",
		b"11111101011011010001010110",
		b"11111101011001001010000101",
		b"11111101010111001001001101",
		b"11111101010101001110110000",
		b"11111101010011011010110011",
		b"11111101010001101101011000",
		b"11111101010000000110100010",
		b"11111101001110100110010100",
		b"11111101001101001100101111",
		b"11111101001011111001110111",
		b"11111101001010101101101100",
		b"11111101001001101000010000",
		b"11111101001000101001100101",
		b"11111101000111110001101011",
		b"11111101000111000000100100",
		b"11111101000110010110001111",
		b"11111101000101110010101101",
		b"11111101000101010101111111",
		b"11111101000101000000000011",
		b"11111101000100110000111010",
		b"11111101000100101000100011",
		b"11111101000100100110111101",
		b"11111101000100101100000110",
		b"11111101000100110111111110",
		b"11111101000101001010100010",
		b"11111101000101100011110001",
		b"11111101000110000011101001",
		b"11111101000110101010001000",
		b"11111101000111010111001010",
		b"11111101001000001010101101",
		b"11111101001001000100101110",
		b"11111101001010000101001010",
		b"11111101001011001011111100",
		b"11111101001100011001000011",
		b"11111101001101101100011001",
		b"11111101001111000101111011",
		b"11111101010000100101100011",
		b"11111101010010001011001111",
		b"11111101010011110110111000",
		b"11111101010101101000011010",
		b"11111101010111011111110000",
		b"11111101011001011100110100",
		b"11111101011011011111100001",
		b"11111101011101100111110010",
		b"11111101011111110101100000",
		b"11111101100010001000100101",
		b"11111101100100100000111010",
		b"11111101100110111110011011",
		b"11111101101001100000111111",
		b"11111101101100001000100001",
		b"11111101101110110100111000",
		b"11111101110001100101111111",
		b"11111101110100011011101110",
		b"11111101110111010101111110",
		b"11111101111010010100100110",
		b"11111101111101010111100001",
		b"11111110000000011110100100",
		b"11111110000011101001101010",
		b"11111110000110111000101001",
		b"11111110001010001011011010",
		b"11111110001101100001110100",
		b"11111110010000111011101111",
		b"11111110010100011001000010",
		b"11111110010111111001100110",
		b"11111110011011011101010001",
		b"11111110011111000011111010",
		b"11111110100010101101011001",
		b"11111110100110011001100101",
		b"11111110101010001000010100",
		b"11111110101101111001011111",
		b"11111110110001101100111011",
		b"11111110110101100010011111",
		b"11111110111001011010000011",
		b"11111110111101010011011101",
		b"11111111000001001110100011",
		b"11111111000101001011001101",
		b"11111111001001001001010001",
		b"11111111001101001000100110",
		b"11111111010001001001000010",
		b"11111111010101001010011011",
		b"11111111011001001100101001",
		b"11111111011101001111100010",
		b"11111111100001010010111101",
		b"11111111100101010110110000",
		b"11111111101001011010110001",
		b"11111111101101011110111000",
		b"11111111110001100010111010",
		b"11111111110101100110110000",
		b"11111111111001101010001110",
		b"11111111111101101101001101",
		b"00000000000001101111100011",
		b"00000000000101110001000110",
		b"00000000001001110001101110",
		b"00000000001101110001010001",
		b"00000000010001101111100111",
		b"00000000010101101100100110",
		b"00000000011001101000000110",
		b"00000000011101100001111110",
		b"00000000100001011010000101",
		b"00000000100101010000010011",
		b"00000000101001000100011111",
		b"00000000101100110110100001",
		b"00000000110000100110010000",
		b"00000000110100010011100101",
		b"00000000110111111110010110",
		b"00000000111011100110011101",
		b"00000000111111001011110001",
		b"00000001000010101110001011",
		b"00000001000110001101100010",
		b"00000001001001101001110000",
		b"00000001001101000010101110",
		b"00000001010000011000010011",
		b"00000001010011101010011000",
		b"00000001010110111000111000",
		b"00000001011010000011101011",
		b"00000001011101001010101010",
		b"00000001100000001101110000",
		b"00000001100011001100110101",
		b"00000001100110000111110100",
		b"00000001101000111110100110",
		b"00000001101011110001000110",
		b"00000001101110011111001111",
		b"00000001110001001000111010",
		b"00000001110011101110000010",
		b"00000001110110001110100011",
		b"00000001111000101010010111",
		b"00000001111011000001011001",
		b"00000001111101010011100110",
		b"00000001111111100000111000",
		b"00000010000001101001001011",
		b"00000010000011101100011101",
		b"00000010000101101010100111",
		b"00000010000111100011101000",
		b"00000010001001010111011011",
		b"00000010001011000101111110",
		b"00000010001100101111001100",
		b"00000010001110010011000101",
		b"00000010001111110001100100",
		b"00000010010001001010101000",
		b"00000010010010011110001110",
		b"00000010010011101100010100",
		b"00000010010100110100111001",
		b"00000010010101110111111010",
		b"00000010010110110101010111",
		b"00000010010111101101001101",
		b"00000010011000011111011101",
		b"00000010011001001100000110",
		b"00000010011001110011000110",
		b"00000010011010010100011110",
		b"00000010011010110000001100",
		b"00000010011011000110010010",
		b"00000010011011010110110000",
		b"00000010011011100001100101",
		b"00000010011011100110110011",
		b"00000010011011100110011010",
		b"00000010011011100000011011",
		b"00000010011011010100111000",
		b"00000010011011000011110010",
		b"00000010011010101101001010",
		b"00000010011010010001000011",
		b"00000010011001101111011110",
		b"00000010011001001000011110",
		b"00000010011000011100000101",
		b"00000010010111101010010101",
		b"00000010010110110011010010",
		b"00000010010101110110111101",
		b"00000010010100110101011011",
		b"00000010010011101110101111",
		b"00000010010010100010111100",
		b"00000010010001010010000101",
		b"00000010001111111100001111",
		b"00000010001110100001011110",
		b"00000010001101000001110101",
		b"00000010001011011101011001",
		b"00000010001001110100001110",
		b"00000010001000000110011010",
		b"00000010000110010100000001",
		b"00000010000100011101000111",
		b"00000010000010100001110010",
		b"00000010000000100010000111",
		b"00000001111110011110001100",
		b"00000001111100010110000101",
		b"00000001111010001001111010",
		b"00000001110111111001101110",
		b"00000001110101100101101001",
		b"00000001110011001101110000",
		b"00000001110000110010001010",
		b"00000001101110010010111100",
		b"00000001101011110000001110",
		b"00000001101001001010000101",
		b"00000001100110100000101000",
		b"00000001100011110011111110",
		b"00000001100001000100001101",
		b"00000001011110010001011101",
		b"00000001011011011011110100",
		b"00000001011000100011011010",
		b"00000001010101101000010110",
		b"00000001010010101010101110",
		b"00000001001111101010101010",
		b"00000001001100101000010001",
		b"00000001001001100011101100",
		b"00000001000110011101000000",
		b"00000001000011010100010111",
		b"00000001000000001001110110",
		b"00000000111100111101100111",
		b"00000000111001101111110000",
		b"00000000110110100000011010",
		b"00000000110011001111101011",
		b"00000000101111111101101100",
		b"00000000101100101010100101",
		b"00000000101001010110011100",
		b"00000000100110000001011011",
		b"00000000100010101011101001",
		b"00000000011111010101001101",
		b"00000000011011111110010000",
		b"00000000011000100110111010",
		b"00000000010101001111010001",
		b"00000000010001110111011110",
		b"00000000001110011111101001",
		b"00000000001011000111111010",
		b"00000000000111110000010111",
		b"00000000000100011001001010",
		b"00000000000001000010011001",
		b"11111111111101101100001100",
		b"11111111111010010110101011",
		b"11111111110111000001111101",
		b"11111111110011101110001010",
		b"11111111110000011011011010",
		b"11111111101101001001110011",
		b"11111111101001111001011100",
		b"11111111100110101010011111",
		b"11111111100011011101000000",
		b"11111111100000010001001000",
		b"11111111011101000110111101",
		b"11111111011001111110100111",
		b"11111111010110111000001100",
		b"11111111010011110011110100",
		b"11111111010000110001100100",
		b"11111111001101110001100011",
		b"11111111001010110011111001",
		b"11111111000111111000101010",
		b"11111111000100111111111111",
		b"11111111000010001001111011",
		b"11111110111111010110100111",
		b"11111110111100100110000111",
		b"11111110111001111000100010",
		b"11111110110111001101111101",
		b"11111110110100100110011110",
		b"11111110110010000010001010",
		b"11111110101111100001000111",
		b"11111110101101000011011001",
		b"11111110101010101001000111",
		b"11111110101000010010010100",
		b"11111110100101111111000101",
		b"11111110100011101111100000",
		b"11111110100001100011101001",
		b"11111110011111011011100011",
		b"11111110011101010111010100",
		b"11111110011011010110111111",
		b"11111110011001011010101000",
		b"11111110010111100010010100",
		b"11111110010101101110000100",
		b"11111110010011111101111110",
		b"11111110010010010010000100",
		b"11111110010000101010011001",
		b"11111110001111000111000000",
		b"11111110001101100111111101",
		b"11111110001100001101010001",
		b"11111110001010110111000000",
		b"11111110001001100101001011",
		b"11111110001000010111110100",
		b"11111110000111001110111110",
		b"11111110000110001010101011",
		b"11111110000101001010111011",
		b"11111110000100001111110001",
		b"11111110000011011001001110",
		b"11111110000010100111010010",
		b"11111110000001111010000000",
		b"11111110000001010001010111",
		b"11111110000000101101011000",
		b"11111110000000001110000100",
		b"11111101111111110011011011",
		b"11111101111111011101011101",
		b"11111101111111001100001010",
		b"11111101111110111111100010",
		b"11111101111110110111100100",
		b"11111101111110110100010000",
		b"11111101111110110101100101",
		b"11111101111110111011100010",
		b"11111101111111000110000111",
		b"11111101111111010101010001",
		b"11111101111111101001000000",
		b"11111110000000000001010011",
		b"11111110000000011110000110",
		b"11111110000000111111011001",
		b"11111110000001100101001010",
		b"11111110000010001111010101",
		b"11111110000010111101111010",
		b"11111110000011110000110110",
		b"11111110000100101000000101",
		b"11111110000101100011100101",
		b"11111110000110100011010100",
		b"11111110000111100111001110",
		b"11111110001000101111010000",
		b"11111110001001111011010110",
		b"11111110001011001011011110",
		b"11111110001100011111100100",
		b"11111110001101110111100011",
		b"11111110001111010011011000",
		b"11111110010000110011000000",
		b"11111110010010010110010101",
		b"11111110010011111101010100",
		b"11111110010101100111111000",
		b"11111110010111010101111101",
		b"11111110011001000111011110",
		b"11111110011010111100010111",
		b"11111110011100110100100010",
		b"11111110011110101111111100",
		b"11111110100000101110011110",
		b"11111110100010110000000100",
		b"11111110100100110100101000",
		b"11111110100110111100000110",
		b"11111110101001000110010111",
		b"11111110101011010011010111",
		b"11111110101101100010111111",
		b"11111110101111110101001011",
		b"11111110110010001001110100",
		b"11111110110100100000110101",
		b"11111110110110111010001000",
		b"11111110111001010101100111",
		b"11111110111011110011001011",
		b"11111110111110010010110000",
		b"11111111000000110100001110",
		b"11111111000011010111100001",
		b"11111111000101111100100000",
		b"11111111001000100011000111",
		b"11111111001011001011001111",
		b"11111111001101110100110010",
		b"11111111010000011111101001",
		b"11111111010011001011101110",
		b"11111111010101111000111011",
		b"11111111011000100111001000",
		b"11111111011011010110010001",
		b"11111111011110000110001110",
		b"11111111100000110110111001",
		b"11111111100011101000001011",
		b"11111111100110011001111110",
		b"11111111101001001100001100",
		b"11111111101011111110101110",
		b"11111111101110110001011101",
		b"11111111110001100100010011",
		b"11111111110100010111001010",
		b"11111111110111001001111011",
		b"11111111111001111100100000",
		b"11111111111100101110110010",
		b"11111111111111100000101100",
		b"00000000000010010010000111",
		b"00000000000101000010111100",
		b"00000000000111110011000101",
		b"00000000001010100010011100",
		b"00000000001101010000111100",
		b"00000000001111111110011101",
		b"00000000010010101010111011",
		b"00000000010101010110001110",
		b"00000000011000000000010001",
		b"00000000011010101000111110",
		b"00000000011101010000001111",
		b"00000000011111110101111111",
		b"00000000100010011010001000",
		b"00000000100100111100100100",
		b"00000000100111011101001110",
		b"00000000101001111100000000",
		b"00000000101100011000110101",
		b"00000000101110110011101000",
		b"00000000110001001100010100",
		b"00000000110011100010110011",
		b"00000000110101110111000000",
		b"00000000111000001000110111",
		b"00000000111010011000010010",
		b"00000000111100100101001110",
		b"00000000111110101111100101",
		b"00000001000000110111010100",
		b"00000001000010111100010101",
		b"00000001000100111110100100",
		b"00000001000110111101111101",
		b"00000001001000111010011101",
		b"00000001001010110011111110",
		b"00000001001100101010011110",
		b"00000001001110011101111001",
		b"00000001010000001110001011",
		b"00000001010001111011010001",
		b"00000001010011100101000111",
		b"00000001010101001011101010",
		b"00000001010110101110110111",
		b"00000001011000001110101011",
		b"00000001011001101011000100",
		b"00000001011011000011111110",
		b"00000001011100011001010111",
		b"00000001011101101011001101",
		b"00000001011110111001011110",
		b"00000001100000000100000111",
		b"00000001100001001011000110",
		b"00000001100010001110011001",
		b"00000001100011001101111111",
		b"00000001100100001001110110",
		b"00000001100101000001111100",
		b"00000001100101110110010001",
		b"00000001100110100110110011",
		b"00000001100111010011100001",
		b"00000001100111111100011010",
		b"00000001101000100001011101",
		b"00000001101001000010101010",
		b"00000001101001100000000001",
		b"00000001101001111001100000",
		b"00000001101010001111001000",
		b"00000001101010100000111001",
		b"00000001101010101110110010",
		b"00000001101010111000110101",
		b"00000001101010111111000000",
		b"00000001101011000001010110",
		b"00000001101010111111110101",
		b"00000001101010111010100000",
		b"00000001101010110001010111",
		b"00000001101010100100011011",
		b"00000001101010010011101110",
		b"00000001101001111111010000",
		b"00000001101001100111000010",
		b"00000001101001001011001000",
		b"00000001101000101011100001",
		b"00000001101000001000010001",
		b"00000001100111100001011000",
		b"00000001100110110110111010",
		b"00000001100110001000110111",
		b"00000001100101010111010011",
		b"00000001100100100010010000",
		b"00000001100011101001110001",
		b"00000001100010101101111000",
		b"00000001100001101110100111",
		b"00000001100000101100000010",
		b"00000001011111100110001101",
		b"00000001011110011101001000",
		b"00000001011101010000111010",
		b"00000001011100000001100011",
		b"00000001011010101111001000",
		b"00000001011001011001101101",
		b"00000001011000000001010100",
		b"00000001010110100110000011",
		b"00000001010101000111111011",
		b"00000001010011100111000010",
		b"00000001010010000011011100",
		b"00000001010000011101001011",
		b"00000001001110110100010110",
		b"00000001001101001000111111",
		b"00000001001011011011001011",
		b"00000001001001101010111111",
		b"00000001000111111000011110",
		b"00000001000110000011101110",
		b"00000001000100001100110011",
		b"00000001000010010011110010",
		b"00000001000000011000110000",
		b"00000000111110011011110000",
		b"00000000111100011100111001",
		b"00000000111010011100001110",
		b"00000000111000011001110110",
		b"00000000110110010101110100",
		b"00000000110100010000001110",
		b"00000000110010001001001010",
		b"00000000110000000000101011",
		b"00000000101101110110110111",
		b"00000000101011101011110100",
		b"00000000101001011111100111",
		b"00000000100111010010010100",
		b"00000000100101000100000010",
		b"00000000100010110100110101",
		b"00000000100000100100110010",
		b"00000000011110010100000000",
		b"00000000011100000010100011",
		b"00000000011001110000100001",
		b"00000000010111011101111110",
		b"00000000010101001011000001",
		b"00000000010010110111101111",
		b"00000000010000100100001100",
		b"00000000001110010000011111",
		b"00000000001011111100101100",
		b"00000000001001101000111010",
		b"00000000000111010101001101",
		b"00000000000101000001101010",
		b"00000000000010101110010111",
		b"00000000000000011011011001",
		b"11111111111110001000110101",
		b"11111111111011110110110000",
		b"11111111111001100101010000",
		b"11111111110111010100011010",
		b"11111111110101000100010010",
		b"11111111110010110100111110",
		b"11111111110000100110100010",
		b"11111111101110011001000100",
		b"11111111101100001100101001",
		b"11111111101010000001010101",
		b"11111111100111110111001101",
		b"11111111100101101110010101",
		b"11111111100011100110110011",
		b"11111111100001100000101100",
		b"11111111011111011100000010",
		b"11111111011101011000111100",
		b"11111111011011010111011110",
		b"11111111011001010111101011",
		b"11111111010111011001101000",
		b"11111111010101011101011010",
		b"11111111010011100011000011",
		b"11111111010001101010101001",
		b"11111111001111110100010000",
		b"11111111001101111111111011",
		b"11111111001100001101101101",
		b"11111111001010011101101100",
		b"11111111001000101111111001",
		b"11111111000111000100011001",
		b"11111111000101011011010000",
		b"11111111000011110100100000",
		b"11111111000010010000001100",
		b"11111111000000101110011001",
		b"11111110111111001111001000",
		b"11111110111101110010011110",
		b"11111110111100011000011100",
		b"11111110111011000001000101",
		b"11111110111001101100011100",
		b"11111110111000011010100100",
		b"11111110110111001011011111",
		b"11111110110101111111001111",
		b"11111110110100110101110110",
		b"11111110110011101111010111",
		b"11111110110010101011110011",
		b"11111110110001101011001101",
		b"11111110110000101101100110",
		b"11111110101111110011000000",
		b"11111110101110111011011100",
		b"11111110101110000110111011",
		b"11111110101101010101100000",
		b"11111110101100100111001011",
		b"11111110101011111011111101",
		b"11111110101011010011111000",
		b"11111110101010101110111100",
		b"11111110101010001101001001",
		b"11111110101001101110100001",
		b"11111110101001010011000100",
		b"11111110101000111010110010",
		b"11111110101000100101101100",
		b"11111110101000010011110001",
		b"11111110101000000101000010",
		b"11111110100111111001100000",
		b"11111110100111110001001000",
		b"11111110100111101011111100",
		b"11111110100111101001111011",
		b"11111110100111101011000100",
		b"11111110100111101111010111",
		b"11111110100111110110110010",
		b"11111110101000000001010110",
		b"11111110101000001111000001",
		b"11111110101000011111110010",
		b"11111110101000110011101000",
		b"11111110101001001010100001",
		b"11111110101001100100011100",
		b"11111110101010000001011001",
		b"11111110101010100001010100",
		b"11111110101011000100001101",
		b"11111110101011101010000001",
		b"11111110101100010010101111",
		b"11111110101100111110010100",
		b"11111110101101101100110000",
		b"11111110101110011101111110",
		b"11111110101111010001111110",
		b"11111110110000001000101100",
		b"11111110110001000010000110",
		b"11111110110001111110001011",
		b"11111110110010111100110110",
		b"11111110110011111110000101",
		b"11111110110101000001110110",
		b"11111110110110001000000110",
		b"11111110110111010000110001",
		b"11111110111000011011110101",
		b"11111110111001101001001110",
		b"11111110111010111000111001",
		b"11111110111100001010110100",
		b"11111110111101011110111010",
		b"11111110111110110101001000",
		b"11111111000000001101011010",
		b"11111111000001100111101110",
		b"11111111000011000100000000",
		b"11111111000100100010001011",
		b"11111111000110000010001100",
		b"11111111000111100100000000",
		b"11111111001001000111100010",
		b"11111111001010101100101111",
		b"11111111001100010011100010",
		b"11111111001101111011111001",
		b"11111111001111100101101101",
		b"11111111010001010000111101",
		b"11111111010010111101100011",
		b"11111111010100101011011100",
		b"11111111010110011010100010",
		b"11111111011000001010110011",
		b"11111111011001111100001010",
		b"11111111011011101110100010",
		b"11111111011101100001110111",
		b"11111111011111010110000110",
		b"11111111100001001011001001",
		b"11111111100011000000111100",
		b"11111111100100110111011100",
		b"11111111100110101110100010",
		b"11111111101000100110001101",
		b"11111111101010011110010110",
		b"11111111101100010110111001",
		b"11111111101110001111110010",
		b"11111111110000001000111110",
		b"11111111110010000010010110",
		b"11111111110011111011111000",
		b"11111111110101110101011110",
		b"11111111110111101111000100",
		b"11111111111001101000100110",
		b"11111111111011100010000000",
		b"11111111111101011011001100",
		b"11111111111111010100001000",
		b"00000000000001001100101111",
		b"00000000000011000100111100",
		b"00000000000100111100101011",
		b"00000000000110110011111000",
		b"00000000001000101010011111",
		b"00000000001010100000011100",
		b"00000000001100010101101010",
		b"00000000001110001010000110",
		b"00000000001111111101101100",
		b"00000000010001110000010111",
		b"00000000010011100010000100",
		b"00000000010101010010101111",
		b"00000000010111000010010100",
		b"00000000011000110000101111",
		b"00000000011010011101111101",
		b"00000000011100001001111001",
		b"00000000011101110100100001",
		b"00000000011111011101110001",
		b"00000000100001000101100100",
		b"00000000100010101011111001",
		b"00000000100100010000101011",
		b"00000000100101110011110110",
		b"00000000100111010101011001",
		b"00000000101000110101010000",
		b"00000000101010010011010111",
		b"00000000101011101111101100",
		b"00000000101101001010001011",
		b"00000000101110100010110010",
		b"00000000101111111001011110",
		b"00000000110001001110001100",
		b"00000000110010100000111010",
		b"00000000110011110001100100",
		b"00000000110101000000001010",
		b"00000000110110001100100111",
		b"00000000110111010110111010",
		b"00000000111000011111000001",
		b"00000000111001100100111001",
		b"00000000111010101000100000",
		b"00000000111011101001110101",
		b"00000000111100101000110101",
		b"00000000111101100101011111",
		b"00000000111110011111110001",
		b"00000000111111010111101001",
		b"00000001000000001101000110",
		b"00000001000001000000000110",
		b"00000001000001110000101000",
		b"00000001000010011110101011",
		b"00000001000011001010001110",
		b"00000001000011110011001111",
		b"00000001000100011001101101",
		b"00000001000100111101101001",
		b"00000001000101011111000000",
		b"00000001000101111101110010",
		b"00000001000110011001111111",
		b"00000001000110110011100110",
		b"00000001000111001010100110",
		b"00000001000111011111000000",
		b"00000001000111110000110011",
		b"00000001000111111111111111",
		b"00000001001000001100100011",
		b"00000001001000010110100001",
		b"00000001001000011101111000",
		b"00000001001000100010101000",
		b"00000001001000100100110010",
		b"00000001001000100100010110",
		b"00000001001000100001010101",
		b"00000001001000011011101110",
		b"00000001001000010011100100",
		b"00000001001000001000110111",
		b"00000001000111111011100111",
		b"00000001000111101011110110",
		b"00000001000111011001100100",
		b"00000001000111000100110011",
		b"00000001000110101101100100",
		b"00000001000110010011111000",
		b"00000001000101110111110001",
		b"00000001000101011001010000",
		b"00000001000100111000010111",
		b"00000001000100010101000111",
		b"00000001000011101111100011",
		b"00000001000011000111101011",
		b"00000001000010011101100001",
		b"00000001000001110001001001",
		b"00000001000001000010100011",
		b"00000001000000010001110001",
		b"00000000111111011110110111",
		b"00000000111110101001110110",
		b"00000000111101110010110000",
		b"00000000111100111001101000",
		b"00000000111011111110100000",
		b"00000000111011000001011011",
		b"00000000111010000010011100",
		b"00000000111001000001100100",
		b"00000000110111111110110111",
		b"00000000110110111010010111",
		b"00000000110101110100000111",
		b"00000000110100101100001010",
		b"00000000110011100010100100",
		b"00000000110010010111010101",
		b"00000000110001001010100011",
		b"00000000101111111100010000",
		b"00000000101110101100011110",
		b"00000000101101011011010001",
		b"00000000101100001000101101",
		b"00000000101010110100110100",
		b"00000000101001011111101010",
		b"00000000101000001001010010",
		b"00000000100110110001101111",
		b"00000000100101011001000101",
		b"00000000100011111111010110",
		b"00000000100010100100100111",
		b"00000000100001001000111011",
		b"00000000011111101100010101",
		b"00000000011110001110111001",
		b"00000000011100110000101011",
		b"00000000011011010001101101",
		b"00000000011001110010000011",
		b"00000000011000010001110001",
		b"00000000010110110000111011",
		b"00000000010101001111100011",
		b"00000000010011101101101111",
		b"00000000010010001011100000",
		b"00000000010000101000111011",
		b"00000000001111000110000011",
		b"00000000001101100010111100",
		b"00000000001011111111101001",
		b"00000000001010011100001111",
		b"00000000001000111000110000",
		b"00000000000111010101010000",
		b"00000000000101110001110010",
		b"00000000000100001110011011",
		b"00000000000010101011001110",
		b"00000000000001001000001110",
		b"11111111111111100101011111",
		b"11111111111110000011000100",
		b"11111111111100100001000000",
		b"11111111111010111111011000",
		b"11111111111001011110001110",
		b"11111111110111111101100101",
		b"11111111110110011101100010",
		b"11111111110100111110001000",
		b"11111111110011011111011001",
		b"11111111110010000001011001",
		b"11111111110000100100001011",
		b"11111111101111000111110010",
		b"11111111101101101100010010",
		b"11111111101100010001101110",
		b"11111111101010111000001000",
		b"11111111101001011111100100",
		b"11111111101000001000000100",
		b"11111111100110110001101100",
		b"11111111100101011100011110",
		b"11111111100100001000011101",
		b"11111111100010110101101100",
		b"11111111100001100100001101",
		b"11111111100000010100000100",
		b"11111111011111000101010010",
		b"11111111011101110111111011",
		b"11111111011100101100000001",
		b"11111111011011100001100110",
		b"11111111011010011000101100",
		b"11111111011001010001010110",
		b"11111111011000001011100111",
		b"11111111010111000111011111",
		b"11111111010110000101000010",
		b"11111111010101000100010010",
		b"11111111010100000101010000",
		b"11111111010011000111111110",
		b"11111111010010001100011110",
		b"11111111010001010010110010",
		b"11111111010000011010111100",
		b"11111111001111100100111101",
		b"11111111001110110000110110",
		b"11111111001101111110101010",
		b"11111111001101001110011010",
		b"11111111001100100000000110",
		b"11111111001011110011110001",
		b"11111111001011001001011011",
		b"11111111001010100001000110",
		b"11111111001001111010110010",
		b"11111111001001010110100001",
		b"11111111001000110100010011",
		b"11111111001000010100001001",
		b"11111111000111110110000101",
		b"11111111000111011010000110",
		b"11111111000111000000001101",
		b"11111111000110101000011011",
		b"11111111000110010010110000",
		b"11111111000101111111001100",
		b"11111111000101101101110001",
		b"11111111000101011110011101",
		b"11111111000101010001010001",
		b"11111111000101000110001110",
		b"11111111000100111101010010",
		b"11111111000100110110011111",
		b"11111111000100110001110011",
		b"11111111000100101111001111",
		b"11111111000100101110110010",
		b"11111111000100110000011100",
		b"11111111000100110100001100",
		b"11111111000100111010000010",
		b"11111111000101000001111101",
		b"11111111000101001011111101",
		b"11111111000101011000000001",
		b"11111111000101100110000111",
		b"11111111000101110110001111",
		b"11111111000110001000011000",
		b"11111111000110011100100001",
		b"11111111000110110010101001",
		b"11111111000111001010101111",
		b"11111111000111100100110000",
		b"11111111001000000000101101",
		b"11111111001000011110100100",
		b"11111111001000111110010011",
		b"11111111001001011111111000",
		b"11111111001010000011010011",
		b"11111111001010101000100001",
		b"11111111001011001111100001",
		b"11111111001011111000010010",
		b"11111111001100100010110000",
		b"11111111001101001110111011",
		b"11111111001101111100110001",
		b"11111111001110101100001111",
		b"11111111001111011101010100",
		b"11111111010000001111111101",
		b"11111111010001000100001001",
		b"11111111010001111001110100",
		b"11111111010010110000111110",
		b"11111111010011101001100100",
		b"11111111010100100011100011",
		b"11111111010101011110111001",
		b"11111111010110011011100100",
		b"11111111010111011001100001",
		b"11111111011000011000101110",
		b"11111111011001011001001001",
		b"11111111011010011010101110",
		b"11111111011011011101011100",
		b"11111111011100100001001111",
		b"11111111011101100110000101",
		b"11111111011110101011111100",
		b"11111111011111110010110000",
		b"11111111100000111010011111",
		b"11111111100010000011000111",
		b"11111111100011001100100100",
		b"11111111100100010110110011",
		b"11111111100101100001110011",
		b"11111111100110101101011111",
		b"11111111100111111001110110",
		b"11111111101001000110110101",
		b"11111111101010010100011000",
		b"11111111101011100010011100",
		b"11111111101100110000111111",
		b"11111111101101111111111111",
		b"11111111101111001111010111",
		b"11111111110000011111000101",
		b"11111111110001101111000111",
		b"11111111110010111111011001",
		b"11111111110100001111111000",
		b"11111111110101100000100010",
		b"11111111110110110001010100",
		b"11111111111000000010001010",
		b"11111111111001010011000010",
		b"11111111111010100011111001",
		b"11111111111011110100101100",
		b"11111111111101000101011000",
		b"11111111111110010101111011",
		b"11111111111111100110010001",
		b"00000000000000110110011000",
		b"00000000000010000110001101",
		b"00000000000011010101101110",
		b"00000000000100100100110110",
		b"00000000000101110011100100",
		b"00000000000111000001110101",
		b"00000000001000001111100111",
		b"00000000001001011100110110",
		b"00000000001010101001100000",
		b"00000000001011110101100010",
		b"00000000001101000000111011",
		b"00000000001110001011100110",
		b"00000000001111010101100010",
		b"00000000010000011110101101",
		b"00000000010001100111000011",
		b"00000000010010101110100011",
		b"00000000010011110101001010",
		b"00000000010100111010110101",
		b"00000000010101111111100011",
		b"00000000010111000011010010",
		b"00000000011000000101111110",
		b"00000000011001000111100110",
		b"00000000011010001000001000",
		b"00000000011011000111100010",
		b"00000000011100000101110001",
		b"00000000011101000010110100",
		b"00000000011101111110101000",
		b"00000000011110111001001101",
		b"00000000011111110010100000",
		b"00000000100000101010011111",
		b"00000000100001100001001000",
		b"00000000100010010110011011",
		b"00000000100011001010010101",
		b"00000000100011111100110100",
		b"00000000100100101101111000",
		b"00000000100101011101011110",
		b"00000000100110001011100110",
		b"00000000100110111000001110",
		b"00000000100111100011010101",
		b"00000000101000001100111001",
		b"00000000101000110100111010",
		b"00000000101001011011010110",
		b"00000000101010000000001101",
		b"00000000101010100011011100",
		b"00000000101011000101000100",
		b"00000000101011100101000100",
		b"00000000101100000011011010",
		b"00000000101100100000000111",
		b"00000000101100111011001000",
		b"00000000101101010100011110",
		b"00000000101101101100001001",
		b"00000000101110000010000111",
		b"00000000101110010110011000",
		b"00000000101110101000111100",
		b"00000000101110111001110010",
		b"00000000101111001000111011",
		b"00000000101111010110010110",
		b"00000000101111100010000011",
		b"00000000101111101100000010",
		b"00000000101111110100010011",
		b"00000000101111111010110101",
		b"00000000101111111111101010",
		b"00000000110000000010110001",
		b"00000000110000000100001011",
		b"00000000110000000011110111",
		b"00000000110000000001110111",
		b"00000000101111111110001010",
		b"00000000101111111000110001",
		b"00000000101111110001101101",
		b"00000000101111101000111110",
		b"00000000101111011110100101",
		b"00000000101111010010100011",
		b"00000000101111000100111000",
		b"00000000101110110101100101",
		b"00000000101110100100101100",
		b"00000000101110010010001100",
		b"00000000101101111110000111",
		b"00000000101101101000011110",
		b"00000000101101010001010011",
		b"00000000101100111000100101",
		b"00000000101100011110010111",
		b"00000000101100000010101010",
		b"00000000101011100101011111",
		b"00000000101011000110110111",
		b"00000000101010100110110100",
		b"00000000101010000101010111",
		b"00000000101001100010100001",
		b"00000000101000111110010101",
		b"00000000101000011000110011",
		b"00000000100111110001111110",
		b"00000000100111001001110110",
		b"00000000100110100000011110",
		b"00000000100101110101111000",
		b"00000000100101001010000101",
		b"00000000100100011101000110",
		b"00000000100011101110111111",
		b"00000000100010111111110000",
		b"00000000100010001111011011",
		b"00000000100001011110000011",
		b"00000000100000101011101010",
		b"00000000011111111000010001",
		b"00000000011111000011111010",
		b"00000000011110001110101000",
		b"00000000011101011000011101",
		b"00000000011100100001011010",
		b"00000000011011101001100010",
		b"00000000011010110000110111",
		b"00000000011001110111011100",
		b"00000000011000111101010001",
		b"00000000011000000010011011",
		b"00000000010111000110111010",
		b"00000000010110001010110001",
		b"00000000010101001110000010",
		b"00000000010100010000110001",
		b"00000000010011010010111101",
		b"00000000010010010100101100",
		b"00000000010001010101111101",
		b"00000000010000010110110100",
		b"00000000001111010111010100",
		b"00000000001110010111011110",
		b"00000000001101010111010101",
		b"00000000001100010110111010",
		b"00000000001011010110010010",
		b"00000000001010010101011101",
		b"00000000001001010100011110",
		b"00000000001000010011010111",
		b"00000000000111010010001011",
		b"00000000000110010000111101",
		b"00000000000101001111101110",
		b"00000000000100001110100000",
		b"00000000000011001101010111",
		b"00000000000010001100010100",
		b"00000000000001001011011001",
		b"00000000000000001010101010",
		b"11111111111111001010000111",
		b"11111111111110001001110100",
		b"11111111111101001001110010",
		b"11111111111100001010000101",
		b"11111111111011001010101101",
		b"11111111111010001011101101",
		b"11111111111001001101001000",
		b"11111111111000001110111111",
		b"11111111110111010001010101",
		b"11111111110110010100001011",
		b"11111111110101010111100100",
		b"11111111110100011011100001",
		b"11111111110011100000000110",
		b"11111111110010100101010011",
		b"11111111110001101011001011",
		b"11111111110000110001101111",
		b"11111111101111111001000001",
		b"11111111101111000001000100",
		b"11111111101110001001111001",
		b"11111111101101010011100010",
		b"11111111101100011110000001",
		b"11111111101011101001010111",
		b"11111111101010110101100110",
		b"11111111101010000010101111",
		b"11111111101001010000110101",
		b"11111111101000011111111001",
		b"11111111100111101111111100",
		b"11111111100111000001000000",
		b"11111111100110010011000110",
		b"11111111100101100110010000",
		b"11111111100100111010011111",
		b"11111111100100001111110101",
		b"11111111100011100110010010",
		b"11111111100010111101111000",
		b"11111111100010010110101000",
		b"11111111100001110000100011",
		b"11111111100001001011101010",
		b"11111111100000100111111111",
		b"11111111100000000101100010",
		b"11111111011111100100010101",
		b"11111111011111000100011000",
		b"11111111011110100101101100",
		b"11111111011110001000010010",
		b"11111111011101101100001010",
		b"11111111011101010001010110",
		b"11111111011100110111110110",
		b"11111111011100011111101011",
		b"11111111011100001000110101",
		b"11111111011011110011010100",
		b"11111111011011011111001010",
		b"11111111011011001100010111",
		b"11111111011010111010111011",
		b"11111111011010101010110110",
		b"11111111011010011100001000",
		b"11111111011010001110110011",
		b"11111111011010000010110110",
		b"11111111011001111000010001",
		b"11111111011001101111000100",
		b"11111111011001100111001111",
		b"11111111011001100000110011",
		b"11111111011001011011101111",
		b"11111111011001011000000011",
		b"11111111011001010101101111",
		b"11111111011001010100110011",
		b"11111111011001010101001110",
		b"11111111011001010111000000",
		b"11111111011001011010001001",
		b"11111111011001011110101001",
		b"11111111011001100100011110",
		b"11111111011001101011101001",
		b"11111111011001110100001001",
		b"11111111011001111101111101",
		b"11111111011010001001000101",
		b"11111111011010010101100000",
		b"11111111011010100011001101",
		b"11111111011010110010001100",
		b"11111111011011000010011011",
		b"11111111011011010011111011",
		b"11111111011011100110101001",
		b"11111111011011111010100110",
		b"11111111011100001111101111",
		b"11111111011100100110000101",
		b"11111111011100111101100110",
		b"11111111011101010110010000",
		b"11111111011101110000000100",
		b"11111111011110001010111111",
		b"11111111011110100111000001",
		b"11111111011111000100001000",
		b"11111111011111100010010100",
		b"11111111100000000001100010",
		b"11111111100000100001110001",
		b"11111111100001000011000000",
		b"11111111100001100101001110",
		b"11111111100010001000011010",
		b"11111111100010101100100001",
		b"11111111100011010001100010",
		b"11111111100011110111011100",
		b"11111111100100011110001110",
		b"11111111100101000101110101",
		b"11111111100101101110010000",
		b"11111111100110010111011110",
		b"11111111100111000001011101",
		b"11111111100111101100001011",
		b"11111111101000010111100111",
		b"11111111101001000011101111",
		b"11111111101001110000100000",
		b"11111111101010011101111011",
		b"11111111101011001011111100",
		b"11111111101011111010100010",
		b"11111111101100101001101011",
		b"11111111101101011001010110",
		b"11111111101110001001100001",
		b"11111111101110111010001001",
		b"11111111101111101011001101",
		b"11111111110000011100101100",
		b"11111111110001001110100011",
		b"11111111110010000000110000",
		b"11111111110010110011010010",
		b"11111111110011100110000111",
		b"11111111110100011001001101",
		b"11111111110101001100100010",
		b"11111111110110000000000101",
		b"11111111110110110011110010",
		b"11111111110111100111101010",
		b"11111111111000011011101000",
		b"11111111111001001111101101",
		b"11111111111010000011110110",
		b"11111111111010111000000001",
		b"11111111111011101100001100",
		b"11111111111100100000010101",
		b"11111111111101010100011011",
		b"11111111111110001000011100",
		b"11111111111110111100010110",
		b"11111111111111110000000111",
		b"00000000000000100011101101",
		b"00000000000001010111000111",
		b"00000000000010001010010010",
		b"00000000000010111101001110",
		b"00000000000011101111111000",
		b"00000000000100100010001111",
		b"00000000000101010100010000",
		b"00000000000110000101111011",
		b"00000000000110110111001101",
		b"00000000000111101000000101",
		b"00000000001000011000100001",
		b"00000000001001001000100000",
		b"00000000001001111000000000",
		b"00000000001010100110111111",
		b"00000000001011010101011100",
		b"00000000001100000011010110",
		b"00000000001100110000101010",
		b"00000000001101011101011000",
		b"00000000001110001001011110",
		b"00000000001110110100111011",
		b"00000000001111011111101100",
		b"00000000010000001001110010",
		b"00000000010000110011001010",
		b"00000000010001011011110011",
		b"00000000010010000011101100",
		b"00000000010010101010110100",
		b"00000000010011010001001001",
		b"00000000010011110110101011",
		b"00000000010100011011011000",
		b"00000000010100111111001110",
		b"00000000010101100010001110",
		b"00000000010110000100010110",
		b"00000000010110100101100101",
		b"00000000010111000101111001",
		b"00000000010111100101010011",
		b"00000000011000000011110001",
		b"00000000011000100001010010",
		b"00000000011000111101110101",
		b"00000000011001011001011010",
		b"00000000011001110100000000",
		b"00000000011010001101100110",
		b"00000000011010100110001100",
		b"00000000011010111101110000",
		b"00000000011011010100010011",
		b"00000000011011101001110011",
		b"00000000011011111110010000",
		b"00000000011100010001101010",
		b"00000000011100100100000001",
		b"00000000011100110101010011",
		b"00000000011101000101100000",
		b"00000000011101010100101001",
		b"00000000011101100010101100",
		b"00000000011101101111101010",
		b"00000000011101111011100010",
		b"00000000011110000110010101",
		b"00000000011110010000000001",
		b"00000000011110011000100111",
		b"00000000011110100000000111",
		b"00000000011110100110100001",
		b"00000000011110101011110101",
		b"00000000011110110000000011",
		b"00000000011110110011001011",
		b"00000000011110110101001100",
		b"00000000011110110110001001",
		b"00000000011110110101111111",
		b"00000000011110110100110001",
		b"00000000011110110010011101",
		b"00000000011110101111000101",
		b"00000000011110101010101001",
		b"00000000011110100101001001",
		b"00000000011110011110100101",
		b"00000000011110010110111110",
		b"00000000011110001110010101",
		b"00000000011110000100101010",
		b"00000000011101111001111110",
		b"00000000011101101110010001",
		b"00000000011101100001100011",
		b"00000000011101010011110110",
		b"00000000011101000101001011",
		b"00000000011100110101100001",
		b"00000000011100100100111011",
		b"00000000011100010011010111",
		b"00000000011100000000111000",
		b"00000000011011101101011111",
		b"00000000011011011001001011",
		b"00000000011011000011111111",
		b"00000000011010101101111010",
		b"00000000011010010110111111",
		b"00000000011001111111001101",
		b"00000000011001100110100111",
		b"00000000011001001101001100",
		b"00000000011000110010111110",
		b"00000000011000010111111111",
		b"00000000010111111100001111",
		b"00000000010111011111110000",
		b"00000000010111000010100010",
		b"00000000010110100100100111",
		b"00000000010110000110000000",
		b"00000000010101100110101110",
		b"00000000010101000110110011",
		b"00000000010100100110010000",
		b"00000000010100000101000101",
		b"00000000010011100011010101",
		b"00000000010011000001000001",
		b"00000000010010011110001010",
		b"00000000010001111010110001",
		b"00000000010001010110111000",
		b"00000000010000110010100000",
		b"00000000010000001101101010",
		b"00000000001111101000011001",
		b"00000000001111000010101100",
		b"00000000001110011100100110",
		b"00000000001101110110001001",
		b"00000000001101001111010101",
		b"00000000001100101000001100",
		b"00000000001100000000101111",
		b"00000000001011011001000001",
		b"00000000001010110001000010",
		b"00000000001010001000110011",
		b"00000000001001100000010111",
		b"00000000001000110111101111",
		b"00000000001000001110111100",
		b"00000000000111100101111111",
		b"00000000000110111100111011",
		b"00000000000110010011110001",
		b"00000000000101101010100001",
		b"00000000000101000001001110",
		b"00000000000100010111111010",
		b"00000000000011101110100100",
		b"00000000000011000101010000",
		b"00000000000010011011111110",
		b"00000000000001110010110000",
		b"00000000000001001001100111",
		b"00000000000000100000100100",
		b"11111111111111110111101010",
		b"11111111111111001110111010",
		b"11111111111110100110010100",
		b"11111111111101111101111010",
		b"11111111111101010101101111",
		b"11111111111100101101110010",
		b"11111111111100000110000101",
		b"11111111111011011110101011",
		b"11111111111010110111100011",
		b"11111111111010010000110000",
		b"11111111111001101010010010",
		b"11111111111001000100001011",
		b"11111111111000011110011100",
		b"11111111110111111001000111",
		b"11111111110111010100001100",
		b"11111111110110101111101101",
		b"11111111110110001011101011",
		b"11111111110101101000000111",
		b"11111111110101000101000010",
		b"11111111110100100010011110",
		b"11111111110100000000011011",
		b"11111111110011011110111011",
		b"11111111110010111101111110",
		b"11111111110010011101100110",
		b"11111111110001111101110011",
		b"11111111110001011110101000",
		b"11111111110001000000000011",
		b"11111111110000100010000111",
		b"11111111110000000100110101",
		b"11111111101111101000001101",
		b"11111111101111001100010000",
		b"11111111101110110000111111",
		b"11111111101110010110011011",
		b"11111111101101111100100100",
		b"11111111101101100011011011",
		b"11111111101101001011000010",
		b"11111111101100110011011000",
		b"11111111101100011100011110",
		b"11111111101100000110010101",
		b"11111111101011110000111110",
		b"11111111101011011100011001",
		b"11111111101011001000100111",
		b"11111111101010110101100111",
		b"11111111101010100011011100",
		b"11111111101010010010000100",
		b"11111111101010000001100001",
		b"11111111101001110001110011",
		b"11111111101001100010111010",
		b"11111111101001010100110111",
		b"11111111101001000111101001",
		b"11111111101000111011010010",
		b"11111111101000101111110001",
		b"11111111101000100101000111",
		b"11111111101000011011010011",
		b"11111111101000010010010110",
		b"11111111101000001010010001",
		b"11111111101000000011000010",
		b"11111111100111111100101011",
		b"11111111100111110111001011",
		b"11111111100111110010100010",
		b"11111111100111101110110000",
		b"11111111100111101011110101",
		b"11111111100111101001110010",
		b"11111111100111101000100101",
		b"11111111100111101000001110",
		b"11111111100111101000101111",
		b"11111111100111101010000101",
		b"11111111100111101100010010",
		b"11111111100111101111010100",
		b"11111111100111110011001100",
		b"11111111100111110111111001",
		b"11111111100111111101011011",
		b"11111111101000000011110001",
		b"11111111101000001010111011",
		b"11111111101000010010111001",
		b"11111111101000011011101010",
		b"11111111101000100101001101",
		b"11111111101000101111100010",
		b"11111111101000111010101001",
		b"11111111101001000110100001",
		b"11111111101001010011001010",
		b"11111111101001100000100010",
		b"11111111101001101110101001",
		b"11111111101001111101011110",
		b"11111111101010001101000010",
		b"11111111101010011101010010",
		b"11111111101010101110001111",
		b"11111111101010111111110111",
		b"11111111101011010010001010",
		b"11111111101011100101000111",
		b"11111111101011111000101101",
		b"11111111101100001100111100",
		b"11111111101100100001110010",
		b"11111111101100110111001110",
		b"11111111101101001101010001",
		b"11111111101101100011111000",
		b"11111111101101111011000011",
		b"11111111101110010010110001",
		b"11111111101110101011000001",
		b"11111111101111000011110010",
		b"11111111101111011101000011",
		b"11111111101111110110110011",
		b"11111111110000010001000001",
		b"11111111110000101011101100",
		b"11111111110001000110110011",
		b"11111111110001100010010101",
		b"11111111110001111110010001",
		b"11111111110010011010100101",
		b"11111111110010110111010001",
		b"11111111110011010100010100",
		b"11111111110011110001101100",
		b"11111111110100001111011001",
		b"11111111110100101101011001",
		b"11111111110101001011101011",
		b"11111111110101101010001111",
		b"11111111110110001001000010",
		b"11111111110110101000000100",
		b"11111111110111000111010011",
		b"11111111110111100110110000",
		b"11111111111000000110010111",
		b"11111111111000100110001001",
		b"11111111111001000110000100",
		b"11111111111001100110000110",
		b"11111111111010000110010000",
		b"11111111111010100110011111",
		b"11111111111011000110110011",
		b"11111111111011100111001010",
		b"11111111111100000111100011",
		b"11111111111100100111111101",
		b"11111111111101001000011000",
		b"11111111111101101000110001",
		b"11111111111110001001001000",
		b"11111111111110101001011011",
		b"11111111111111001001101010",
		b"11111111111111101001110011",
		b"00000000000000001001110101",
		b"00000000000000101001110000",
		b"00000000000001001001100001",
		b"00000000000001101001001001",
		b"00000000000010001000100101",
		b"00000000000010100111110110",
		b"00000000000011000110111001",
		b"00000000000011100101101110",
		b"00000000000100000100010100",
		b"00000000000100100010101001",
		b"00000000000101000000101101",
		b"00000000000101011110100000",
		b"00000000000101111011111110",
		b"00000000000110011001001001",
		b"00000000000110110101111111",
		b"00000000000111010010011111",
		b"00000000000111101110100111",
		b"00000000001000001010011000",
		b"00000000001000100101110001",
		b"00000000001001000000101111",
		b"00000000001001011011010100",
		b"00000000001001110101011101",
		b"00000000001010001111001010",
		b"00000000001010101000011010",
		b"00000000001011000001001101",
		b"00000000001011011001100001",
		b"00000000001011110001010111",
		b"00000000001100001000101100",
		b"00000000001100011111100001",
		b"00000000001100110101110101",
		b"00000000001101001011100111",
		b"00000000001101100000110110",
		b"00000000001101110101100011",
		b"00000000001110001001101100",
		b"00000000001110011101010000",
		b"00000000001110110000010000",
		b"00000000001111000010101011",
		b"00000000001111010100100000",
		b"00000000001111100101101110",
		b"00000000001111110110010110",
		b"00000000010000000110010111",
		b"00000000010000010101110000",
		b"00000000010000100100100001",
		b"00000000010000110010101010",
		b"00000000010001000000001011",
		b"00000000010001001101000010",
		b"00000000010001011001010000",
		b"00000000010001100100110101",
		b"00000000010001101111101111",
		b"00000000010001111010000000",
		b"00000000010010000011100111",
		b"00000000010010001100100011",
		b"00000000010010010100110101",
		b"00000000010010011100011100",
		b"00000000010010100011011000",
		b"00000000010010101001101001",
		b"00000000010010101111010000",
		b"00000000010010110100001011",
		b"00000000010010111000011100",
		b"00000000010010111100000010",
		b"00000000010010111110111101",
		b"00000000010011000001001101",
		b"00000000010011000010110010",
		b"00000000010011000011101101",
		b"00000000010011000011111101",
		b"00000000010011000011100011",
		b"00000000010011000010011111",
		b"00000000010011000000110000",
		b"00000000010010111110011000",
		b"00000000010010111011010111",
		b"00000000010010110111101100",
		b"00000000010010110011011000",
		b"00000000010010101110011011",
		b"00000000010010101000110111",
		b"00000000010010100010101010",
		b"00000000010010011011110101",
		b"00000000010010010100011001",
		b"00000000010010001100010111",
		b"00000000010010000011101110",
		b"00000000010001111010011111",
		b"00000000010001110000101011",
		b"00000000010001100110010001",
		b"00000000010001011011010011",
		b"00000000010001001111110001",
		b"00000000010001000011101100",
		b"00000000010000110111000100",
		b"00000000010000101001111001",
		b"00000000010000011100001101",
		b"00000000010000001101111111",
		b"00000000001111111111010001",
		b"00000000001111110000000011",
		b"00000000001111100000010110",
		b"00000000001111010000001010",
		b"00000000001110111111100000",
		b"00000000001110101110011010",
		b"00000000001110011100110110",
		b"00000000001110001010110111",
		b"00000000001101111000011101",
		b"00000000001101100101101000",
		b"00000000001101010010011010",
		b"00000000001100111110110011",
		b"00000000001100101010110101",
		b"00000000001100010110011110",
		b"00000000001100000001110010",
		b"00000000001011101100110000",
		b"00000000001011010111011001",
		b"00000000001011000001101110",
		b"00000000001010101011110000",
		b"00000000001010010101011111",
		b"00000000001001111110111101",
		b"00000000001001101000001010",
		b"00000000001001010001001000",
		b"00000000001000111001110110",
		b"00000000001000100010010111",
		b"00000000001000001010101010",
		b"00000000000111110010110001",
		b"00000000000111011010101101",
		b"00000000000111000010011101",
		b"00000000000110101010000101",
		b"00000000000110010001100011",
		b"00000000000101111000111010",
		b"00000000000101100000001001",
		b"00000000000101000111010010",
		b"00000000000100101110010110",
		b"00000000000100010101010110",
		b"00000000000011111100010010",
		b"00000000000011100011001011",
		b"00000000000011001010000011",
		b"00000000000010110000111001",
		b"00000000000010010111110000",
		b"00000000000001111110101000",
		b"00000000000001100101100001",
		b"00000000000001001100011101",
		b"00000000000000110011011100",
		b"00000000000000011010100000",
		b"00000000000000000001101001",
		b"11111111111111101000111000",
		b"11111111111111010000001110",
		b"11111111111110110111101011",
		b"11111111111110011111010001",
		b"11111111111110000111000000",
		b"11111111111101101110111001",
		b"11111111111101010110111101",
		b"11111111111100111111001101",
		b"11111111111100100111101001",
		b"11111111111100010000010010",
		b"11111111111011111001001010",
		b"11111111111011100010010000",
		b"11111111111011001011100101",
		b"11111111111010110101001011",
		b"11111111111010011111000001",
		b"11111111111010001001001001",
		b"11111111111001110011100100",
		b"11111111111001011110010001",
		b"11111111111001001001010010",
		b"11111111111000110100101000",
		b"11111111111000100000010010",
		b"11111111111000001100010001",
		b"11111111110111111000100111",
		b"11111111110111100101010100",
		b"11111111110111010010011000",
		b"11111111110110111111110011",
		b"11111111110110101101100111",
		b"11111111110110011011110100",
		b"11111111110110001010011011",
		b"11111111110101111001011011",
		b"11111111110101101000110110",
		b"11111111110101011000101100",
		b"11111111110101001000111101",
		b"11111111110100111001101011",
		b"11111111110100101010110100",
		b"11111111110100011100011010",
		b"11111111110100001110011101",
		b"11111111110100000000111101",
		b"11111111110011110011111011",
		b"11111111110011100111010111",
		b"11111111110011011011010010",
		b"11111111110011001111101011",
		b"11111111110011000100100011",
		b"11111111110010111001111011",
		b"11111111110010101111110010",
		b"11111111110010100110001000",
		b"11111111110010011100111111",
		b"11111111110010010100010110",
		b"11111111110010001100001100",
		b"11111111110010000100100100",
		b"11111111110001111101011100",
		b"11111111110001110110110100",
		b"11111111110001110000101110",
		b"11111111110001101011001000",
		b"11111111110001100110000011",
		b"11111111110001100001100000",
		b"11111111110001011101011101",
		b"11111111110001011001111011",
		b"11111111110001010110111010",
		b"11111111110001010100011011",
		b"11111111110001010010011100",
		b"11111111110001010000111110",
		b"11111111110001010000000001",
		b"11111111110001001111100101",
		b"11111111110001001111101001",
		b"11111111110001010000001101",
		b"11111111110001010001010010",
		b"11111111110001010010111000",
		b"11111111110001010100111101",
		b"11111111110001010111100010",
		b"11111111110001011010100110",
		b"11111111110001011110001010",
		b"11111111110001100010001101",
		b"11111111110001100110101111",
		b"11111111110001101011101111",
		b"11111111110001110001001101",
		b"11111111110001110111001010",
		b"11111111110001111101100100",
		b"11111111110010000100011011",
		b"11111111110010001011110000",
		b"11111111110010010011100001",
		b"11111111110010011011101110",
		b"11111111110010100100010111",
		b"11111111110010101101011011",
		b"11111111110010110110111010",
		b"11111111110011000000110100",
		b"11111111110011001011001000",
		b"11111111110011010101110110",
		b"11111111110011100000111100",
		b"11111111110011101100011100",
		b"11111111110011111000010011",
		b"11111111110100000100100010",
		b"11111111110100010001001001",
		b"11111111110100011110000110",
		b"11111111110100101011011001",
		b"11111111110100111001000010",
		b"11111111110101000111000000",
		b"11111111110101010101010010",
		b"11111111110101100011111000",
		b"11111111110101110010110001",
		b"11111111110110000001111101",
		b"11111111110110010001011100",
		b"11111111110110100001001011",
		b"11111111110110110001001100",
		b"11111111110111000001011101",
		b"11111111110111010001111101",
		b"11111111110111100010101101",
		b"11111111110111110011101011",
		b"11111111111000000100110111",
		b"11111111111000010110010000",
		b"11111111111000100111110101",
		b"11111111111000111001100110",
		b"11111111111001001011100010",
		b"11111111111001011101101001",
		b"11111111111001101111111001",
		b"11111111111010000010010011",
		b"11111111111010010100110101",
		b"11111111111010100111011111",
		b"11111111111010111010010000",
		b"11111111111011001101001000",
		b"11111111111011100000000101",
		b"11111111111011110011001000",
		b"11111111111100000110001111",
		b"11111111111100011001011010",
		b"11111111111100101100101000",
		b"11111111111100111111111000",
		b"11111111111101010011001010",
		b"11111111111101100110011101",
		b"11111111111101111001110001",
		b"11111111111110001101000100",
		b"11111111111110100000010110",
		b"11111111111110110011100111",
		b"11111111111111000110110110",
		b"11111111111111011010000010",
		b"11111111111111101101001010",
		b"00000000000000000000001110",
		b"00000000000000010011001101",
		b"00000000000000100110000111",
		b"00000000000000111000111011",
		b"00000000000001001011101000",
		b"00000000000001011110001110",
		b"00000000000001110000101100",
		b"00000000000010000011000010",
		b"00000000000010010101001110",
		b"00000000000010100111010001",
		b"00000000000010111001001001",
		b"00000000000011001010110111",
		b"00000000000011011100011001",
		b"00000000000011101101110000",
		b"00000000000011111110111010",
		b"00000000000100001111110110",
		b"00000000000100100000100110",
		b"00000000000100110001000111",
		b"00000000000101000001011001",
		b"00000000000101010001011101",
		b"00000000000101100001010001",
		b"00000000000101110000110100",
		b"00000000000110000000001000",
		b"00000000000110001111001010",
		b"00000000000110011101111011",
		b"00000000000110101100011010",
		b"00000000000110111010100111",
		b"00000000000111001000100001",
		b"00000000000111010110001000",
		b"00000000000111100011011011",
		b"00000000000111110000011011",
		b"00000000000111111101000110",
		b"00000000001000001001011101",
		b"00000000001000010101011111",
		b"00000000001000100001001011",
		b"00000000001000101100100010",
		b"00000000001000110111100011",
		b"00000000001001000010001110",
		b"00000000001001001100100011",
		b"00000000001001010110100000",
		b"00000000001001100000000111",
		b"00000000001001101001010111",
		b"00000000001001110010001111",
		b"00000000001001111010110000",
		b"00000000001010000010111001",
		b"00000000001010001010101001",
		b"00000000001010010010000010",
		b"00000000001010011001000010",
		b"00000000001010011111101010",
		b"00000000001010100101111010",
		b"00000000001010101011110000",
		b"00000000001010110001001110",
		b"00000000001010110110010011",
		b"00000000001010111010111111",
		b"00000000001010111111010010",
		b"00000000001011000011001100",
		b"00000000001011000110101100",
		b"00000000001011001001110100",
		b"00000000001011001100100010",
		b"00000000001011001110111000",
		b"00000000001011010000110100",
		b"00000000001011010010010111",
		b"00000000001011010011100001",
		b"00000000001011010100010011",
		b"00000000001011010100101011",
		b"00000000001011010100101011",
		b"00000000001011010100010001",
		b"00000000001011010011100000",
		b"00000000001011010010010110",
		b"00000000001011010000110011",
		b"00000000001011001110111001",
		b"00000000001011001100100110",
		b"00000000001011001001111011",
		b"00000000001011000110111001",
		b"00000000001011000011100000",
		b"00000000001010111111101111",
		b"00000000001010111011100111",
		b"00000000001010110111001001",
		b"00000000001010110010010100",
		b"00000000001010101101001001",
		b"00000000001010100111100111",
		b"00000000001010100001110000",
		b"00000000001010011011100100",
		b"00000000001010010101000010",
		b"00000000001010001110001100",
		b"00000000001010000111000001",
		b"00000000001001111111100001",
		b"00000000001001110111101110",
		b"00000000001001101111101000",
		b"00000000001001100111001110",
		b"00000000001001011110100010",
		b"00000000001001010101100011",
		b"00000000001001001100010010",
		b"00000000001001000010101111",
		b"00000000001000111000111100",
		b"00000000001000101110110111",
		b"00000000001000100100100010",
		b"00000000001000011001111101",
		b"00000000001000001111001000",
		b"00000000001000000100000100",
		b"00000000000111111000110010",
		b"00000000000111101101010001",
		b"00000000000111100001100010",
		b"00000000000111010101100110",
		b"00000000000111001001011101",
		b"00000000000110111101001000",
		b"00000000000110110000100110",
		b"00000000000110100011111001",
		b"00000000000110010111000001",
		b"00000000000110001001111111",
		b"00000000000101111100110010",
		b"00000000000101101111011100",
		b"00000000000101100001111101",
		b"00000000000101010100010101",
		b"00000000000101000110100110",
		b"00000000000100111000101110",
		b"00000000000100101010110000",
		b"00000000000100011100101010",
		b"00000000000100001110011111",
		b"00000000000100000000001111",
		b"00000000000011110001111001",
		b"00000000000011100011011110",
		b"00000000000011010101000000",
		b"00000000000011000110011110",
		b"00000000000010110111111001",
		b"00000000000010101001010010",
		b"00000000000010011010101000",
		b"00000000000010001011111101",
		b"00000000000001111101010001",
		b"00000000000001101110100101",
		b"00000000000001011111111000",
		b"00000000000001010001001100",
		b"00000000000001000010100001",
		b"00000000000000110011111000",
		b"00000000000000100101010000",
		b"00000000000000010110101011",
		b"00000000000000001000001001",
		b"11111111111111111001101010",
		b"11111111111111101011001111",
		b"11111111111111011100111001",
		b"11111111111111001110100111",
		b"11111111111111000000011011",
		b"11111111111110110010010100",
		b"11111111111110100100010100",
		b"11111111111110010110011010",
		b"11111111111110001000101000",
		b"11111111111101111010111101",
		b"11111111111101101101011010",
		b"11111111111101011111111111",
		b"11111111111101010010101110",
		b"11111111111101000101100101",
		b"11111111111100111000100110",
		b"11111111111100101011110010",
		b"11111111111100011111000111",
		b"11111111111100010010101000",
		b"11111111111100000110010011",
		b"11111111111011111010001011",
		b"11111111111011101110001110",
		b"11111111111011100010011101",
		b"11111111111011010110111010",
		b"11111111111011001011100011",
		b"11111111111011000000011001",
		b"11111111111010110101011101",
		b"11111111111010101010110000",
		b"11111111111010100000010000",
		b"11111111111010010101111111",
		b"11111111111010001011111101",
		b"11111111111010000010001001",
		b"11111111111001111000100110",
		b"11111111111001101111010010",
		b"11111111111001100110001110",
		b"11111111111001011101011010",
		b"11111111111001010100110110",
		b"11111111111001001100100011",
		b"11111111111001000100100001",
		b"11111111111000111100101111",
		b"11111111111000110101001111",
		b"11111111111000101110000001",
		b"11111111111000100111000100",
		b"11111111111000100000011001",
		b"11111111111000011001111111",
		b"11111111111000010011111000",
		b"11111111111000001110000011",
		b"11111111111000001000100000",
		b"11111111111000000011001111",
		b"11111111110111111110010001",
		b"11111111110111111001100101",
		b"11111111110111110101001101",
		b"11111111110111110001000111",
		b"11111111110111101101010011",
		b"11111111110111101001110011",
		b"11111111110111100110100101",
		b"11111111110111100011101011",
		b"11111111110111100001000011",
		b"11111111110111011110101111",
		b"11111111110111011100101101",
		b"11111111110111011010111110",
		b"11111111110111011001100010",
		b"11111111110111011000011001",
		b"11111111110111010111100011",
		b"11111111110111010111000000",
		b"11111111110111010110110000",
		b"11111111110111010110110010",
		b"11111111110111010111000111",
		b"11111111110111010111101110",
		b"11111111110111011000101000",
		b"11111111110111011001110100",
		b"11111111110111011011010011",
		b"11111111110111011101000011",
		b"11111111110111011111000110",
		b"11111111110111100001011010",
		b"11111111110111100100000000",
		b"11111111110111100110110111",
		b"11111111110111101010000000",
		b"11111111110111101101011010",
		b"11111111110111110001000101",
		b"11111111110111110101000000",
		b"11111111110111111001001101",
		b"11111111110111111101101001",
		b"11111111111000000010010110",
		b"11111111111000000111010011",
		b"11111111111000001100100000",
		b"11111111111000010001111100",
		b"11111111111000010111100111",
		b"11111111111000011101100001",
		b"11111111111000100011101010",
		b"11111111111000101010000001",
		b"11111111111000110000100111",
		b"11111111111000110111011010",
		b"11111111111000111110011011",
		b"11111111111001000101101010",
		b"11111111111001001101000101",
		b"11111111111001010100101101",
		b"11111111111001011100100010",
		b"11111111111001100100100010",
		b"11111111111001101100101111",
		b"11111111111001110101000111",
		b"11111111111001111101101010",
		b"11111111111010000110011000",
		b"11111111111010001111010000",
		b"11111111111010011000010010",
		b"11111111111010100001011111",
		b"11111111111010101010110100",
		b"11111111111010110100010011",
		b"11111111111010111101111011",
		b"11111111111011000111101011",
		b"11111111111011010001100011",
		b"11111111111011011011100010",
		b"11111111111011100101101001",
		b"11111111111011101111110111",
		b"11111111111011111010001100",
		b"11111111111100000100100110",
		b"11111111111100001111000111",
		b"11111111111100011001101100",
		b"11111111111100100100010111",
		b"11111111111100101111000111",
		b"11111111111100111001111011",
		b"11111111111101000100110011",
		b"11111111111101001111101110",
		b"11111111111101011010101101",
		b"11111111111101100101101110",
		b"11111111111101110000110010",
		b"11111111111101111011111000",
		b"11111111111110000110111111",
		b"11111111111110010010001000",
		b"11111111111110011101010010",
		b"11111111111110101000011100",
		b"11111111111110110011100110",
		b"11111111111110111110110000",
		b"11111111111111001001111010",
		b"11111111111111010101000010",
		b"11111111111111100000001010",
		b"11111111111111101011001111",
		b"11111111111111110110010011",
		b"00000000000000000001010100",
		b"00000000000000001100010010",
		b"00000000000000010111001101",
		b"00000000000000100010000101",
		b"00000000000000101100111001",
		b"00000000000000110111101001",
		b"00000000000001000010010100",
		b"00000000000001001100111010",
		b"00000000000001010111011100",
		b"00000000000001100001110111",
		b"00000000000001101100001101",
		b"00000000000001110110011101",
		b"00000000000010000000100110",
		b"00000000000010001010101000",
		b"00000000000010010100100100",
		b"00000000000010011110011000",
		b"00000000000010101000000100",
		b"00000000000010110001101000",
		b"00000000000010111011000100",
		b"00000000000011000100011000",
		b"00000000000011001101100011",
		b"00000000000011010110100100",
		b"00000000000011011111011100",
		b"00000000000011101000001011",
		b"00000000000011110000110000",
		b"00000000000011111001001010",
		b"00000000000100000001011011",
		b"00000000000100001001100000",
		b"00000000000100010001011011",
		b"00000000000100011001001011",
		b"00000000000100100000110000",
		b"00000000000100101000001001",
		b"00000000000100101111010110",
		b"00000000000100110110011000",
		b"00000000000100111101001110",
		b"00000000000101000011110111",
		b"00000000000101001010010100",
		b"00000000000101010000100101",
		b"00000000000101010110101001",
		b"00000000000101011100100000",
		b"00000000000101100010001010",
		b"00000000000101100111100111",
		b"00000000000101101100110110",
		b"00000000000101110001111001",
		b"00000000000101110110101101",
		b"00000000000101111011010100",
		b"00000000000101111111101110",
		b"00000000000110000011111010",
		b"00000000000110000111110111",
		b"00000000000110001011100111",
		b"00000000000110001111001001",
		b"00000000000110010010011101",
		b"00000000000110010101100010",
		b"00000000000110011000011010",
		b"00000000000110011011000011",
		b"00000000000110011101011110",
		b"00000000000110011111101011",
		b"00000000000110100001101001",
		b"00000000000110100011011001",
		b"00000000000110100100111011",
		b"00000000000110100110001110",
		b"00000000000110100111010011",
		b"00000000000110101000001010",
		b"00000000000110101000110011",
		b"00000000000110101001001101",
		b"00000000000110101001011010",
		b"00000000000110101001011000",
		b"00000000000110101001001000",
		b"00000000000110101000101010",
		b"00000000000110100111111110",
		b"00000000000110100111000100",
		b"00000000000110100101111101",
		b"00000000000110100100101000",
		b"00000000000110100011000101",
		b"00000000000110100001010101",
		b"00000000000110011111010111",
		b"00000000000110011101001100",
		b"00000000000110011010110100",
		b"00000000000110011000001111",
		b"00000000000110010101011101",
		b"00000000000110010010011111",
		b"00000000000110001111010011",
		b"00000000000110001011111100",
		b"00000000000110001000011000",
		b"00000000000110000100101000",
		b"00000000000110000000101100",
		b"00000000000101111100100100",
		b"00000000000101111000010000",
		b"00000000000101110011110010",
		b"00000000000101101111000111",
		b"00000000000101101010010010",
		b"00000000000101100101010010",
		b"00000000000101100000001000",
		b"00000000000101011010110011",
		b"00000000000101010101010100",
		b"00000000000101001111101011",
		b"00000000000101001001111000",
		b"00000000000101000011111011",
		b"00000000000100111101110110",
		b"00000000000100110111100111",
		b"00000000000100110001001111",
		b"00000000000100101010101111",
		b"00000000000100100100000110",
		b"00000000000100011101010110",
		b"00000000000100010110011101",
		b"00000000000100001111011101",
		b"00000000000100001000010101",
		b"00000000000100000001000111",
		b"00000000000011111001110001",
		b"00000000000011110010010101",
		b"00000000000011101010110011",
		b"00000000000011100011001011",
		b"00000000000011011011011101",
		b"00000000000011010011101001",
		b"00000000000011001011110000",
		b"00000000000011000011110011",
		b"00000000000010111011110000",
		b"00000000000010110011101001",
		b"00000000000010101011011111",
		b"00000000000010100011010000",
		b"00000000000010011010111110",
		b"00000000000010010010101000",
		b"00000000000010001010010000",
		b"00000000000010000001110100",
		b"00000000000001111001010111",
		b"00000000000001110000110111",
		b"00000000000001101000010110",
		b"00000000000001011111110010",
		b"00000000000001010111001110",
		b"00000000000001001110101000",
		b"00000000000001000110000010",
		b"00000000000000111101011100",
		b"00000000000000110100110101",
		b"00000000000000101100001110",
		b"00000000000000100011101000",
		b"00000000000000011011000010",
		b"00000000000000010010011110",
		b"00000000000000001001111010",
		b"00000000000000000001011000",
		b"11111111111111111000111000",
		b"11111111111111110000011010",
		b"11111111111111100111111110",
		b"11111111111111011111100100",
		b"11111111111111010111001110",
		b"11111111111111001110111010",
		b"11111111111111000110101010",
		b"11111111111110111110011101",
		b"11111111111110110110010100",
		b"11111111111110101110010000",
		b"11111111111110100110001111",
		b"11111111111110011110010011",
		b"11111111111110010110011100",
		b"11111111111110001110101010",
		b"11111111111110000110111101",
		b"11111111111101111111010110",
		b"11111111111101110111110101",
		b"11111111111101110000011001",
		b"11111111111101101001000011",
		b"11111111111101100001110100",
		b"11111111111101011010101100",
		b"11111111111101010011101010",
		b"11111111111101001100101111",
		b"11111111111101000101111100",
		b"11111111111100111111001111",
		b"11111111111100111000101011",
		b"11111111111100110010001110",
		b"11111111111100101011111001",
		b"11111111111100100101101100",
		b"11111111111100011111100111",
		b"11111111111100011001101011",
		b"11111111111100010011110111",
		b"11111111111100001110001101",
		b"11111111111100001000101011",
		b"11111111111100000011010010",
		b"11111111111011111110000010",
		b"11111111111011111000111011",
		b"11111111111011110011111110",
		b"11111111111011101111001011",
		b"11111111111011101010100001",
		b"11111111111011100110000001",
		b"11111111111011100001101011",
		b"11111111111011011101011111",
		b"11111111111011011001011101",
		b"11111111111011010101100110",
		b"11111111111011010001111000",
		b"11111111111011001110010101",
		b"11111111111011001010111101",
		b"11111111111011000111101111",
		b"11111111111011000100101100",
		b"11111111111011000001110011",
		b"11111111111010111111000101",
		b"11111111111010111100100010",
		b"11111111111010111010001001",
		b"11111111111010110111111100",
		b"11111111111010110101111001",
		b"11111111111010110100000010",
		b"11111111111010110010010101",
		b"11111111111010110000110011",
		b"11111111111010101111011100",
		b"11111111111010101110010000",
		b"11111111111010101101001111",
		b"11111111111010101100011001",
		b"11111111111010101011101111",
		b"11111111111010101011001111",
		b"11111111111010101010111010",
		b"11111111111010101010110000",
		b"11111111111010101010110000",
		b"11111111111010101010111100",
		b"11111111111010101011010010",
		b"11111111111010101011110100",
		b"11111111111010101100100000",
		b"11111111111010101101010110",
		b"11111111111010101110010111",
		b"11111111111010101111100011",
		b"11111111111010110000111001",
		b"11111111111010110010011010",
		b"11111111111010110100000101",
		b"11111111111010110101111010",
		b"11111111111010110111111001",
		b"11111111111010111010000011",
		b"11111111111010111100010110",
		b"11111111111010111110110011",
		b"11111111111011000001011010",
		b"11111111111011000100001011",
		b"11111111111011000111000101",
		b"11111111111011001010001001",
		b"11111111111011001101010101",
		b"11111111111011010000101011",
		b"11111111111011010100001010",
		b"11111111111011010111110010",
		b"11111111111011011011100011",
		b"11111111111011011111011100",
		b"11111111111011100011011110",
		b"11111111111011100111101000",
		b"11111111111011101011111010",
		b"11111111111011110000010101",
		b"11111111111011110100110111",
		b"11111111111011111001100001",
		b"11111111111011111110010010",
		b"11111111111100000011001011",
		b"11111111111100001000001011",
		b"11111111111100001101010010",
		b"11111111111100010010100000",
		b"11111111111100010111110101",
		b"11111111111100011101010000",
		b"11111111111100100010110001",
		b"11111111111100101000011000",
		b"11111111111100101110000110",
		b"11111111111100110011111001",
		b"11111111111100111001110010",
		b"11111111111100111111110000",
		b"11111111111101000101110011",
		b"11111111111101001011111100",
		b"11111111111101010010001001",
		b"11111111111101011000011010",
		b"11111111111101011110110000",
		b"11111111111101100101001010",
		b"11111111111101101011101001",
		b"11111111111101110010001010",
		b"11111111111101111000110000",
		b"11111111111101111111011001",
		b"11111111111110000110000101",
		b"11111111111110001100110100",
		b"11111111111110010011100101",
		b"11111111111110011010011001",
		b"11111111111110100001010000",
		b"11111111111110101000001000",
		b"11111111111110101111000011",
		b"11111111111110110101111111",
		b"11111111111110111100111101",
		b"11111111111111000011111100",
		b"11111111111111001010111011",
		b"11111111111111010001111100",
		b"11111111111111011000111110",
		b"11111111111111011111111111",
		b"11111111111111100111000001",
		b"11111111111111101110000011",
		b"11111111111111110101000101",
		b"11111111111111111100000111",
		b"00000000000000000011000111",
		b"00000000000000001010000111",
		b"00000000000000010001000110",
		b"00000000000000011000000100",
		b"00000000000000011111000000",
		b"00000000000000100101111011",
		b"00000000000000101100110100",
		b"00000000000000110011101011",
		b"00000000000000111010011111",
		b"00000000000001000001010001",
		b"00000000000001001000000001",
		b"00000000000001001110101110",
		b"00000000000001010101011000",
		b"00000000000001011011111110",
		b"00000000000001100010100010",
		b"00000000000001101001000001",
		b"00000000000001101111011101",
		b"00000000000001110101110110",
		b"00000000000001111100001010",
		b"00000000000010000010011010",
		b"00000000000010001000100101",
		b"00000000000010001110101100",
		b"00000000000010010100101110",
		b"00000000000010011010101011",
		b"00000000000010100000100100",
		b"00000000000010100110010111",
		b"00000000000010101100000100",
		b"00000000000010110001101101",
		b"00000000000010110111001111",
		b"00000000000010111100101100",
		b"00000000000011000010000010",
		b"00000000000011000111010011",
		b"00000000000011001100011101",
		b"00000000000011010001100001",
		b"00000000000011010110011111",
		b"00000000000011011011010110",
		b"00000000000011100000000110",
		b"00000000000011100100101111",
		b"00000000000011101001010010",
		b"00000000000011101101101101",
		b"00000000000011110010000001",
		b"00000000000011110110001110",
		b"00000000000011111010010011",
		b"00000000000011111110010001",
		b"00000000000100000010000111",
		b"00000000000100000101110110",
		b"00000000000100001001011100",
		b"00000000000100001100111011",
		b"00000000000100010000010010",
		b"00000000000100010011100001",
		b"00000000000100010110101000",
		b"00000000000100011001100111",
		b"00000000000100011100011101",
		b"00000000000100011111001011",
		b"00000000000100100001110001",
		b"00000000000100100100001110",
		b"00000000000100100110100011",
		b"00000000000100101000110000",
		b"00000000000100101010110100",
		b"00000000000100101100101111",
		b"00000000000100101110100001",
		b"00000000000100110000001011",
		b"00000000000100110001101101",
		b"00000000000100110011000101",
		b"00000000000100110100010101",
		b"00000000000100110101011100",
		b"00000000000100110110011011",
		b"00000000000100110111010000",
		b"00000000000100110111111101",
		b"00000000000100111000100001",
		b"00000000000100111000111100",
		b"00000000000100111001001110",
		b"00000000000100111001011000",
		b"00000000000100111001011001",
		b"00000000000100111001010001",
		b"00000000000100111001000000",
		b"00000000000100111000100111",
		b"00000000000100111000000100",
		b"00000000000100110111011010",
		b"00000000000100110110100110",
		b"00000000000100110101101010",
		b"00000000000100110100100110",
		b"00000000000100110011011001",
		b"00000000000100110010000011",
		b"00000000000100110000100101",
		b"00000000000100101110111111",
		b"00000000000100101101010000",
		b"00000000000100101011011001",
		b"00000000000100101001011010",
		b"00000000000100100111010010",
		b"00000000000100100101000011",
		b"00000000000100100010101011",
		b"00000000000100100000001100",
		b"00000000000100011101100101",
		b"00000000000100011010110110",
		b"00000000000100010111111111",
		b"00000000000100010101000001",
		b"00000000000100010001111011",
		b"00000000000100001110101101",
		b"00000000000100001011011001",
		b"00000000000100000111111100",
		b"00000000000100000100011001",
		b"00000000000100000000101111",
		b"00000000000011111100111110",
		b"00000000000011111001000110",
		b"00000000000011110101000111",
		b"00000000000011110001000001",
		b"00000000000011101100110101",
		b"00000000000011101000100010",
		b"00000000000011100100001001",
		b"00000000000011011111101010",
		b"00000000000011011011000101",
		b"00000000000011010110011010",
		b"00000000000011010001101001",
		b"00000000000011001100110010",
		b"00000000000011000111110101",
		b"00000000000011000010110011",
		b"00000000000010111101101100",
		b"00000000000010111000011111",
		b"00000000000010110011001101",
		b"00000000000010101101110111",
		b"00000000000010101000011011",
		b"00000000000010100010111011",
		b"00000000000010011101010110",
		b"00000000000010010111101100",
		b"00000000000010010001111110",
		b"00000000000010001100001100",
		b"00000000000010000110010110",
		b"00000000000010000000011101",
		b"00000000000001111010011111",
		b"00000000000001110100011110",
		b"00000000000001101110011001",
		b"00000000000001101000010000",
		b"00000000000001100010000101",
		b"00000000000001011011110111",
		b"00000000000001010101100101",
		b"00000000000001001111010001",
		b"00000000000001001000111010",
		b"00000000000001000010100001",
		b"00000000000000111100000101",
		b"00000000000000110101100111",
		b"00000000000000101111000111",
		b"00000000000000101000100101",
		b"00000000000000100010000001",
		b"00000000000000011011011011",
		b"00000000000000010100110100",
		b"00000000000000001110001100",
		b"00000000000000000111100011",
		b"00000000000000000000111000",
		b"11111111111111111010001100",
		b"11111111111111110011100000",
		b"11111111111111101100110011",
		b"11111111111111100110000101",
		b"11111111111111011111010111",
		b"11111111111111011000101001",
		b"11111111111111010001111010",
		b"11111111111111001011001100",
		b"11111111111111000100011110",
		b"11111111111110111101110000",
		b"11111111111110110111000010",
		b"11111111111110110000010101",
		b"11111111111110101001101001",
		b"11111111111110100010111110",
		b"11111111111110011100010011",
		b"11111111111110010101101010",
		b"11111111111110001111000010",
		b"11111111111110001000011011",
		b"11111111111110000001110101",
		b"11111111111101111011010010",
		b"11111111111101110100101111",
		b"11111111111101101110001111",
		b"11111111111101100111110001",
		b"11111111111101100001010100",
		b"11111111111101011010111010",
		b"11111111111101010100100010",
		b"11111111111101001110001101",
		b"11111111111101000111111010",
		b"11111111111101000001101010",
		b"11111111111100111011011100",
		b"11111111111100110101010001",
		b"11111111111100101111001010",
		b"11111111111100101001000101",
		b"11111111111100100011000011",
		b"11111111111100011101000101",
		b"11111111111100010111001010",
		b"11111111111100010001010010",
		b"11111111111100001011011110",
		b"11111111111100000101101110",
		b"11111111111100000000000001",
		b"11111111111011111010011000",
		b"11111111111011110100110011",
		b"11111111111011101111010010",
		b"11111111111011101001110101",
		b"11111111111011100100011100",
		b"11111111111011011111001000",
		b"11111111111011011001110111",
		b"11111111111011010100101011",
		b"11111111111011001111100100",
		b"11111111111011001010100001",
		b"11111111111011000101100010",
		b"11111111111011000000101001",
		b"11111111111010111011110011",
		b"11111111111010110111000011",
		b"11111111111010110010011000",
		b"11111111111010101101110001",
		b"11111111111010101001001111",
		b"11111111111010100100110011",
		b"11111111111010100000011011",
		b"11111111111010011100001001",
		b"11111111111010010111111011",
		b"11111111111010010011110011",
		b"11111111111010001111110000",
		b"11111111111010001011110010",
		b"11111111111010000111111010",
		b"11111111111010000100000111",
		b"11111111111010000000011001",
		b"11111111111001111100110001",
		b"11111111111001111001001110",
		b"11111111111001110101110001",
		b"11111111111001110010011001",
		b"11111111111001101111000111",
		b"11111111111001101011111010",
		b"11111111111001101000110011",
		b"11111111111001100101110001",
		b"11111111111001100010110101",
		b"11111111111001011111111111",
		b"11111111111001011101001110",
		b"11111111111001011010100011",
		b"11111111111001010111111101",
		b"11111111111001010101011110",
		b"11111111111001010011000011",
		b"11111111111001010000101111",
		b"11111111111001001110100000",
		b"11111111111001001100010111",
		b"11111111111001001010010011",
		b"11111111111001001000010101",
		b"11111111111001000110011101",
		b"11111111111001000100101010",
		b"11111111111001000010111101",
		b"11111111111001000001010110",
		b"11111111111000111111110100",
		b"11111111111000111110010111",
		b"11111111111000111101000001",
		b"11111111111000111011101111",
		b"11111111111000111010100100",
		b"11111111111000111001011110",
		b"11111111111000111000011101",
		b"11111111111000110111100001",
		b"11111111111000110110101100",
		b"11111111111000110101111011",
		b"11111111111000110101010000",
		b"11111111111000110100101010",
		b"11111111111000110100001001",
		b"11111111111000110011101110",
		b"11111111111000110011011000",
		b"11111111111000110011000111",
		b"11111111111000110010111011",
		b"11111111111000110010110101",
		b"11111111111000110010110011",
		b"11111111111000110010110111",
		b"11111111111000110010111111",
		b"11111111111000110011001100",
		b"11111111111000110011011110",
		b"11111111111000110011110101",
		b"11111111111000110100010001",
		b"11111111111000110100110010",
		b"11111111111000110101010111",
		b"11111111111000110110000001",
		b"11111111111000110110101111",
		b"11111111111000110111100010",
		b"11111111111000111000011010",
		b"11111111111000111001010101",
		b"11111111111000111010010110",
		b"11111111111000111011011010",
		b"11111111111000111100100011",
		b"11111111111000111101110000",
		b"11111111111000111111000001",
		b"11111111111001000000010110",
		b"11111111111001000001101111",
		b"11111111111001000011001100",
		b"11111111111001000100101101",
		b"11111111111001000110010010",
		b"11111111111001000111111010",
		b"11111111111001001001100110",
		b"11111111111001001011010110",
		b"11111111111001001101001010",
		b"11111111111001001111000000",
		b"11111111111001010000111011",
		b"11111111111001010010111000",
		b"11111111111001010100111001",
		b"11111111111001010110111101",
		b"11111111111001011001000101",
		b"11111111111001011011001111",
		b"11111111111001011101011101",
		b"11111111111001011111101101",
		b"11111111111001100010000000",
		b"11111111111001100100010111",
		b"11111111111001100110101111",
		b"11111111111001101001001011",
		b"11111111111001101011101001",
		b"11111111111001101110001010",
		b"11111111111001110000101101",
		b"11111111111001110011010011",
		b"11111111111001110101111011",
		b"11111111111001111000100101",
		b"11111111111001111011010001",
		b"11111111111001111110000000",
		b"11111111111010000000110001",
		b"11111111111010000011100011",
		b"11111111111010000110011000",
		b"11111111111010001001001110",
		b"11111111111010001100000111",
		b"11111111111010001111000001",
		b"11111111111010010001111100",
		b"11111111111010010100111010",
		b"11111111111010010111111000",
		b"11111111111010011010111001",
		b"11111111111010011101111010",
		b"11111111111010100000111101",
		b"11111111111010100100000010",
		b"11111111111010100111000111",
		b"11111111111010101010001110",
		b"11111111111010101101010101",
		b"11111111111010110000011110",
		b"11111111111010110011101000",
		b"11111111111010110110110010",
		b"11111111111010111001111110",
		b"11111111111010111101001010",
		b"11111111111011000000010111",
		b"11111111111011000011100100",
		b"11111111111011000110110010",
		b"11111111111011001010000001",
		b"11111111111011001101010000",
		b"11111111111011010000011111",
		b"11111111111011010011101111",
		b"11111111111011010110111111",
		b"11111111111011011010010000",
		b"11111111111011011101100000",
		b"11111111111011100000110001",
		b"11111111111011100100000010",
		b"11111111111011100111010011",
		b"11111111111011101010100100",
		b"11111111111011101101110100",
		b"11111111111011110001000101",
		b"11111111111011110100010101",
		b"11111111111011110111100101",
		b"11111111111011111010110101",
		b"11111111111011111110000101",
		b"11111111111100000001010100",
		b"11111111111100000100100011",
		b"11111111111100000111110001",
		b"11111111111100001010111111",
		b"11111111111100001110001100",
		b"11111111111100010001011001",
		b"11111111111100010100100101",
		b"11111111111100010111110001",
		b"11111111111100011010111011",
		b"11111111111100011110000101",
		b"11111111111100100001001110",
		b"11111111111100100100010111",
		b"11111111111100100111011110",
		b"11111111111100101010100100",
		b"11111111111100101101101010",
		b"11111111111100110000101111",
		b"11111111111100110011110010",
		b"11111111111100110110110101",
		b"11111111111100111001110110",
		b"11111111111100111100110111",
		b"11111111111100111111110110",
		b"11111111111101000010110100",
		b"11111111111101000101110001",
		b"11111111111101001000101100",
		b"11111111111101001011100111",
		b"11111111111101001110100000",
		b"11111111111101010001010111",
		b"11111111111101010100001110",
		b"11111111111101010111000011",
		b"11111111111101011001110111",
		b"11111111111101011100101001",
		b"11111111111101011111011010",
		b"11111111111101100010001001",
		b"11111111111101100100110111",
		b"11111111111101100111100100",
		b"11111111111101101010001111",
		b"11111111111101101100111000",
		b"11111111111101101111100000",
		b"11111111111101110010000110",
		b"11111111111101110100101011",
		b"11111111111101110111001110",
		b"11111111111101111001110000",
		b"11111111111101111100010000",
		b"11111111111101111110101111",
		b"11111111111110000001001011",
		b"11111111111110000011100110",
		b"11111111111110000110000000",
		b"11111111111110001000011000",
		b"11111111111110001010101110",
		b"11111111111110001101000010",
		b"11111111111110001111010101",
		b"11111111111110010001100110",
		b"11111111111110010011110110",
		b"11111111111110010110000011",
		b"11111111111110011000001111",
		b"11111111111110011010011010",
		b"11111111111110011100100010",
		b"11111111111110011110101001",
		b"11111111111110100000101110",
		b"11111111111110100010110010",
		b"11111111111110100100110011",
		b"11111111111110100110110011",
		b"11111111111110101000110010",
		b"11111111111110101010101110",
		b"11111111111110101100101001",
		b"11111111111110101110100010",
		b"11111111111110110000011001",
		b"11111111111110110010001111",
		b"11111111111110110100000011",
		b"11111111111110110101110101",
		b"11111111111110110111100101",
		b"11111111111110111001010100",
		b"11111111111110111011000001",
		b"11111111111110111100101101",
		b"11111111111110111110010111",
		b"11111111111110111111111111",
		b"11111111111111000001100101",
		b"11111111111111000011001010",
		b"11111111111111000100101101",
		b"11111111111111000110001110",
		b"11111111111111000111101110",
		b"11111111111111001001001100",
		b"11111111111111001010101001",
		b"11111111111111001100000100",
		b"11111111111111001101011101",
		b"11111111111111001110110101",
		b"11111111111111010000001011",
		b"11111111111111010001100000",
		b"11111111111111010010110011",
		b"11111111111111010100000101",
		b"11111111111111010101010101",
		b"11111111111111010110100011",
		b"11111111111111010111110000",
		b"11111111111111011000111100",
		b"11111111111111011010000110",
		b"11111111111111011011001110",
		b"11111111111111011100010101",
		b"11111111111111011101011011",
		b"11111111111111011110011111",
		b"11111111111111011111100010",
		b"11111111111111100000100100",
		b"11111111111111100001100100",
		b"11111111111111100010100011",
		b"11111111111111100011100000",
		b"11111111111111100100011100",
		b"11111111111111100101010111",
		b"11111111111111100110010000",
		b"11111111111111100111001000",
		b"11111111111111100111111111",
		b"11111111111111101000110101",
		b"11111111111111101001101001",
		b"11111111111111101010011100",
		b"11111111111111101011001110",
		b"11111111111111101011111111",
		b"11111111111111101100101111",
		b"11111111111111101101011101",
		b"11111111111111101110001010",
		b"11111111111111101110110110",
		b"11111111111111101111100001",
		b"11111111111111110000001011",
		b"11111111111111110000110100",
		b"11111111111111110001011100",
		b"11111111111111110010000011",
		b"11111111111111110010101000",
		b"11111111111111110011001101",
		b"11111111111111110011110001",
		b"11111111111111110100010011",
		b"11111111111111110100110101",
		b"11111111111111110101010110",
		b"11111111111111110101110110",
		b"11111111111111110110010101",
		b"11111111111111110110110011",
		b"11111111111111110111010000",
		b"11111111111111110111101100",
		b"11111111111111111000001000",
		b"11111111111111111000100010",
		b"11111111111111111000111100",
		b"11111111111111111001010101",
		b"11111111111111111001101101",
		b"11111111111111111010000100",
		b"11111111111111111010011011",
		b"11111111111111111010110001",
		b"11111111111111111011000110",
		b"11111111111111111011011010",
		b"11111111111111111011101110",
		b"11111111111111111100000001",
		b"11111111111111111100010011",
		b"11111111111111111100100101",
		b"11111111111111111100110110",
		b"11111111111111111101000111",
		b"11111111111111111101010111",
		b"11111111111111111101100110",
		b"11111111111111111101110100",
		b"11111111111111111110000010",
		b"11111111111111111110010000",
		b"11111111111111111110011101",
		b"11111111111111111110101001",
		b"11111111111111111110110101",
		b"11111111111111111111000001",
		b"11111111111111111111001100",
		b"11111111111111111111010110",
		b"11111111111111111111100000",
		b"11111111111111111111101001",
		b"11111111111111111111110011",
		b"11111111111111111111111011",
		b"00000000000000000000000011",
		b"00000000000000000000001011",
		b"00000000000000000000010011",
		b"00000000000000000000011010",
		b"00000000000000000000100000",
		b"00000000000000000000100111",
		b"00000000000000000000101100",
		b"00000000000000000000110010",
		b"00000000000000000000110111",
		b"00000000000000000000111100",
		b"00000000000000000001000001",
		b"00000000000000000001000101",
		b"00000000000000000001001001",
		b"00000000000000000001001101",
		b"00000000000000000001010000",
		b"00000000000000000001010100",
		b"00000000000000000001010111",
		b"00000000000000000001011001",
		b"00000000000000000001011100",
		b"00000000000000000001011110",
		b"00000000000000000001100000",
		b"00000000000000000001100010",
		b"00000000000000000001100100",
		b"00000000000000000001100101",
		b"00000000000000000001100110",
		b"00000000000000000001100111",
		b"00000000000000000001101000",
		b"00000000000000000001101001",
		b"00000000000000000001101010",
		b"00000000000000000001101010",
		b"00000000000000000001101010",
		b"00000000000000000001101010",
		b"00000000000000000001101010",
		b"00000000000000000001101010",
		b"00000000000000000001101010",
		b"00000000000000000001101010",
		b"00000000000000000001101001",
		b"00000000000000000001101001",
		b"00000000000000000001101000",
		b"00000000000000000001100111",
		b"00000000000000000001100110",
		b"00000000000000000001100110",
		b"00000000000000000001100101",
		b"00000000000000000001100011",
		b"00000000000000000001100010",
		b"00000000000000000001100001",
		b"00000000000000000001100000",
		b"00000000000000000001011111",
		b"00000000000000000001011101",
		b"00000000000000000001011100",
		b"00000000000000000001011010",
		b"00000000000000000001011001",
		b"00000000000000000001010111",
		b"00000000000000000001010110",
		b"00000000000000000001010100",
		b"00000000000000000001010011",
		b"00000000000000000001010001",
		b"00000000000000000001010000",
		b"00000000000000000001001110",
		b"00000000000000000001001100",
		b"00000000000000000001001011",
		b"00000000000000000001001001",
		b"00000000000000000001000111",
		b"00000000000000000001000110",
		b"00000000000000000001000100",
		b"00000000000000000001000010",
		b"00000000000000000001000000",
		b"00000000000000000000111111",
		b"00000000000000000000111101",
		b"00000000000000000000111011",
		b"00000000000000000000111010",
		b"00000000000000000000111000",
		b"00000000000000000000110110",
		b"00000000000000000000110101",
		b"00000000000000000000110011",
		b"00000000000000000000110010",
		b"00000000000000000000110000",
		b"00000000000000000000101111",
		b"00000000000000000000101101",
		b"00000000000000000000101100",
		b"00000000000000000000101010",
		b"00000000000000000000101001",
		b"00000000000000000000100111",
		b"00000000000000000000100110",
		b"00000000000000000000100100",
		b"00000000000000000000100011",
		b"00000000000000000000100010",
		b"00000000000000000000100000",
		b"00000000000000000000011111",
		b"00000000000000000000011110",
		b"00000000000000000000011100",
		b"00000000000000000000011011",
		b"00000000000000000000011010",
		b"00000000000000000000011001",
		b"00000000000000000000011000",
		b"00000000000000000000010111",
		b"00000000000000000000010110",
		b"00000000000000000000010100",
		b"00000000000000000000010011",
		b"00000000000000000000010010"
	);

end src_rom_pkg;