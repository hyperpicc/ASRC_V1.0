library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package src_rom_pkg is

	constant COE_WIDTH	: integer := 26;
	constant COE_CENTRE	: signed( 25 downto 0 ) := b"01111111010111000010100100";

	type COE_ROM_TYPE is array( 4095 downto 0 ) of signed( 25 downto 0 );
	constant COE_ROM	 : COE_ROM_TYPE := (
		b"01111111010110010001101110",
		b"01111111010011111111010000",
		b"01111111010000001011001100",
		b"01111111001010110101101000",
		b"01111111000011111110101011",
		b"01111110111011100110011110",
		b"01111110110001101101001101",
		b"01111110100110010011000101",
		b"01111110011001011000010111",
		b"01111110001010111101010100",
		b"01111101111011000010010001",
		b"01111101101001100111100011",
		b"01111101010110101101100010",
		b"01111101000010010100101001",
		b"01111100101100011101010011",
		b"01111100010101001000000000",
		b"01111011111100010101001110",
		b"01111011100010000101100001",
		b"01111011000110011001011101",
		b"01111010101001010001100111",
		b"01111010001010101110101001",
		b"01111001101010110001001011",
		b"01111001001001011001111011",
		b"01111000100110101001100101",
		b"01111000000010100000111011",
		b"01110111011101000000101101",
		b"01110110110110001001101111",
		b"01110110001101111100110111",
		b"01110101100100011010111011",
		b"01110100111001100100110101",
		b"01110100001101011011100000",
		b"01110011011111111111111001",
		b"01110010110001010010111011",
		b"01110010000001010101101010",
		b"01110001010000001001000101",
		b"01110000011101101110001111",
		b"01101111101010000110001111",
		b"01101110110101010010001010",
		b"01101101111111010011001000",
		b"01101101001000001010010010",
		b"01101100001111111000110101",
		b"01101011010110011111111011",
		b"01101010011100000000110011",
		b"01101001100000011100101101",
		b"01101000100011110100111001",
		b"01100111100110001010101001",
		b"01100110100111011111010000",
		b"01100101100111110100000100",
		b"01100100100111001010011001",
		b"01100011100101100011100111",
		b"01100010100011000001000111",
		b"01100001011111100100010001",
		b"01100000011011001110100001",
		b"01011111010110000001010001",
		b"01011110001111111101111111",
		b"01011101001001000110000111",
		b"01011100000001011011001010",
		b"01011010111000111110100101",
		b"01011001101111110001111001",
		b"01011000100101110110101000",
		b"01010111011011001110010100",
		b"01010110001111111010011111",
		b"01010101000011111100101101",
		b"01010011110111010110100010",
		b"01010010101010001001100100",
		b"01010001011100010111010111",
		b"01010000001110000001100001",
		b"01001110111111001001101010",
		b"01001101101111110001010111",
		b"01001100011111111010010001",
		b"01001011001111100110000000",
		b"01001001111110110110001100",
		b"01001000101101101100011110",
		b"01000111011100001010011110",
		b"01000110001010010001110110",
		b"01000100111000000100001111",
		b"01000011100101100011010011",
		b"01000010010010110000101011",
		b"01000000111111101110000001",
		b"00111111101100011100111111",
		b"00111110011000111111001111",
		b"00111101000101010110011010",
		b"00111011110001100100001011",
		b"00111010011101101010001010",
		b"00111001001001101010000010",
		b"00110111110101100101011011",
		b"00110110100001011101111111",
		b"00110101001101010101010110",
		b"00110011111001001101001001",
		b"00110010100101000110111111",
		b"00110001010001000100100001",
		b"00101111111101000111010101",
		b"00101110101001010001000011",
		b"00101101010101100011010000",
		b"00101100000001111111100011",
		b"00101010101110100111011111",
		b"00101001011011011100101100",
		b"00101000001000100000101010",
		b"00100110110101110100111110",
		b"00100101100011011011001010",
		b"00100100010001010100101111",
		b"00100010111111100011001111",
		b"00100001101110001000001010",
		b"00100000011101000100111110",
		b"00011111001100011011001010",
		b"00011101111100001100001011",
		b"00011100101100011001011101",
		b"00011011011101000100011011",
		b"00011010001110001110011111",
		b"00011000111111111001000011",
		b"00010111110010000101011110",
		b"00010110100100110101001000",
		b"00010101011000001001010101",
		b"00010100001100000011011011",
		b"00010011000000100100101101",
		b"00010001110101101110011100",
		b"00010000101011100001111010",
		b"00001111100010000000010101",
		b"00001110011001001010111011",
		b"00001101010001000010111010",
		b"00001100001001101001011101",
		b"00001011000010111111101100",
		b"00001001111101000110110010",
		b"00001000110111111111110100",
		b"00000111110011101011111000",
		b"00000110110000001100000010",
		b"00000101101101100001010100",
		b"00000100101011101100101101",
		b"00000011101010101111010011",
		b"00000010101010101001111100",
		b"00000001101011011101100111",
		b"00000000101101001011001110",
		b"11111111101111110011101010",
		b"11111110110011010111110010",
		b"11111101110111111000011011",
		b"11111100111101010110011010",
		b"11111100000011110010011111",
		b"11111011001011001101011100",
		b"11111010010011100111111110",
		b"11111001011101000010110010",
		b"11111000100111011110100100",
		b"11110111110010111011111100",
		b"11110110111111011011100001",
		b"11110110001100111101111010",
		b"11110101011011100011101010",
		b"11110100101011001101010011",
		b"11110011111011111011010110",
		b"11110011001101101110001111",
		b"11110010100000100110011101",
		b"11110001110100100100011001",
		b"11110001001001101000011101",
		b"11110000011111110010111111",
		b"11101111110111000100010101",
		b"11101111001111011100110010",
		b"11101110101000111100100111",
		b"11101110000011100100000011",
		b"11101101011111010011010101",
		b"11101100111100001010101001",
		b"11101100011010001010001000",
		b"11101011111001010001111001",
		b"11101011011001100010001010",
		b"11101010111010111010110101",
		b"11101010011101011100000001",
		b"11101010000001000101110001",
		b"11101001100101111000000001",
		b"11101001001011110010110001",
		b"11101000110010110101111011",
		b"11101000011011000001011010",
		b"11101000000100010101000100",
		b"11100111101110110000110001",
		b"11100111011010010100010100",
		b"11100111000110111111100001",
		b"11100110110100110010001001",
		b"11100110100011101011111010",
		b"11100110010011101100100010",
		b"11100110000100110011101110",
		b"11100101110111000001000111",
		b"11100101101010010100010111",
		b"11100101011110101101000011",
		b"11100101010100001010110010",
		b"11100101001010101101001000",
		b"11100101000010010011100101",
		b"11100100111010111101101100",
		b"11100100110100101010111011",
		b"11100100101111011010110000",
		b"11100100101011001100100111",
		b"11100100100111111111111010",
		b"11100100100101110100000010",
		b"11100100100100101000011000",
		b"11100100100100011100010010",
		b"11100100100101001111000101",
		b"11100100100111000000000001",
		b"11100100101001101110100010",
		b"11100100101101011001101110",
		b"11100100110010000000111001",
		b"11100100110111100011010010",
		b"11100100111110000000000110",
		b"11100101000101010110100001",
		b"11100101001101100101101110",
		b"11100101010110101100110111",
		b"11100101100000101011000011",
		b"11100101101011011111011011",
		b"11100101110111001001000101",
		b"11100110000011100111000111",
		b"11100110010000111000100100",
		b"11100110011110111100100001",
		b"11100110101101110010000000",
		b"11100110111101011000000010",
		b"11100111001101101101101001",
		b"11100111011110110001110100",
		b"11100111110000100011100010",
		b"11101000000011000001110010",
		b"11101000010110001011100010",
		b"11101000101001111111101110",
		b"11101000111110011101010011",
		b"11101001010011100011001100",
		b"11101001101001010000010100",
		b"11101001111111100011100110",
		b"11101010010110011011111011",
		b"11101010101101111000001101",
		b"11101011000101110111010100",
		b"11101011011110011000001010",
		b"11101011110111011001100101",
		b"11101100010000111010011101",
		b"11101100101010111001101110",
		b"11101101000101010110001000",
		b"11101101100000001110100100",
		b"11101101111011100001111010",
		b"11101110010111001110111111",
		b"11101110110011010100101010",
		b"11101111001111110001110001",
		b"11101111101100100101001000",
		b"11110000001001101101100111",
		b"11110000100111001010000010",
		b"11110001000100111001001111",
		b"11110001100010111010000101",
		b"11110010000001001011011001",
		b"11110010011111101100000000",
		b"11110010111110011010110001",
		b"11110011011101010110100010",
		b"11110011111100011110001001",
		b"11110100011011110000011101",
		b"11110100111011001100010100",
		b"11110101011010110000100110",
		b"11110101111010011100001011",
		b"11110110011010001101111001",
		b"11110110111010000100101001",
		b"11110111011001111111010011",
		b"11110111111001111100110001",
		b"11111000011001111011111011",
		b"11111000111001111011101101",
		b"11111001011001111010111111",
		b"11111001111001111000101110",
		b"11111010011001110011110100",
		b"11111010111001101011001110",
		b"11111011011001011101111001",
		b"11111011111001001010110011",
		b"11111100011000110000111000",
		b"11111100111000001111001001",
		b"11111101010111100100100100",
		b"11111101110110110000001011",
		b"11111110010101110000111110",
		b"11111110110100100101111111",
		b"11111111010011001110010001",
		b"11111111110001101000111001",
		b"00000000001111110100111010",
		b"00000000101101110001011001",
		b"00000001001011011101011110",
		b"00000001101000111000010000",
		b"00000010000110000000110110",
		b"00000010100010110110011011",
		b"00000010111111011000001001",
		b"00000011011011100101001010",
		b"00000011110111011100101100",
		b"00000100010010111101111100",
		b"00000100101110001000001000",
		b"00000101001000111010100000",
		b"00000101100011010100010100",
		b"00000101111101010100111000",
		b"00000110010110111011011101",
		b"00000110110000000111011001",
		b"00000111001000110111111111",
		b"00000111100001001100101000",
		b"00000111111001000100101010",
		b"00001000010000011111011111",
		b"00001000100111011100100000",
		b"00001000111101111011001010",
		b"00001001010011111010111001",
		b"00001001101001011011001011",
		b"00001001111110011011100000",
		b"00001010010010111011010111",
		b"00001010100110111010010010",
		b"00001010111010010111110101",
		b"00001011001101010011100011",
		b"00001011011111101101000011",
		b"00001011110001100011111100",
		b"00001100000010110111110101",
		b"00001100010011101000011000",
		b"00001100100011110101010000",
		b"00001100110011011110001010",
		b"00001101000010100010110010",
		b"00001101010001000010111000",
		b"00001101011110111110001100",
		b"00001101101100010100011111",
		b"00001101111001000101100100",
		b"00001110000101010001001111",
		b"00001110010000110111010101",
		b"00001110011011110111101110",
		b"00001110100110010010010001",
		b"00001110110000000110110111",
		b"00001110111001010101011100",
		b"00001111000001111101111011",
		b"00001111001010000000010010",
		b"00001111010001011100011110",
		b"00001111011000010010100000",
		b"00001111011110100010011001",
		b"00001111100100001100001011",
		b"00001111101001001111111010",
		b"00001111101101101101101010",
		b"00001111110001100101100010",
		b"00001111110100110111101001",
		b"00001111110111100100000111",
		b"00001111111001101011000110",
		b"00001111111011001100110001",
		b"00001111111100001001010100",
		b"00001111111100100000111101",
		b"00001111111100010011111001",
		b"00001111111011100010011000",
		b"00001111111010001100101011",
		b"00001111111000010011000100",
		b"00001111110101110101110101",
		b"00001111110010110101010010",
		b"00001111101111010001110001",
		b"00001111101011001011100111",
		b"00001111100110100011001011",
		b"00001111100001011000110110",
		b"00001111011011101101000001",
		b"00001111010101100000000101",
		b"00001111001110110010011110",
		b"00001111000111100100100111",
		b"00001110111111110110111101",
		b"00001110110111101001111111",
		b"00001110101110111110001010",
		b"00001110100101110011111111",
		b"00001110011100001011111101",
		b"00001110010010000110100110",
		b"00001110000111100100011011",
		b"00001101111100100101111111",
		b"00001101110001001011110110",
		b"00001101100101010110100100",
		b"00001101011001000110101101",
		b"00001101001100011100111001",
		b"00001100111111011001101010",
		b"00001100110001111101101011",
		b"00001100100100001001100001",
		b"00001100010101111101110101",
		b"00001100000111011011001111",
		b"00001011111000100010011001",
		b"00001011101001010011111100",
		b"00001011011001110000100011",
		b"00001011001001111000110111",
		b"00001010111001101101100101",
		b"00001010101001001111010111",
		b"00001010011000011110111001",
		b"00001010000111011100111000",
		b"00001001110110001010000001",
		b"00001001100100100111000000",
		b"00001001010010110100100010",
		b"00001001000000110011010101",
		b"00001000101110100100000110",
		b"00001000011100000111100100",
		b"00001000001001011110011101",
		b"00000111110110101001011111",
		b"00000111100011101001011001",
		b"00000111010000011110111000",
		b"00000110111101001010101100",
		b"00000110101001101101100100",
		b"00000110010110001000001110",
		b"00000110000010011011011001",
		b"00000101101110100111110100",
		b"00000101011010101110001110",
		b"00000101000110101111010101",
		b"00000100110010101011111000",
		b"00000100011110100100100110",
		b"00000100001010011010001100",
		b"00000011110110001101011010",
		b"00000011100001111110111110",
		b"00000011001101101111100110",
		b"00000010111001011111111110",
		b"00000010100101010000110101",
		b"00000010010001000010111000",
		b"00000001111100110110110011",
		b"00000001101000101101010100",
		b"00000001010100100111000111",
		b"00000001000000100100110111",
		b"00000000101100100111010000",
		b"00000000011000101110111110",
		b"00000000000100111100101011",
		b"11111111110001010001000001",
		b"11111111011101101100101011",
		b"11111111001010010000010010",
		b"11111110110110111100011111",
		b"11111110100011110001111010",
		b"11111110010000110001001010",
		b"11111101111101111010111001",
		b"11111101101011001111101011",
		b"11111101011000110000001000",
		b"11111101000110011100110101",
		b"11111100110100010110010111",
		b"11111100100010011101010011",
		b"11111100010000110010001011",
		b"11111011111111010101100011",
		b"11111011101110000111111110",
		b"11111011011101001001111110",
		b"11111011001100011100000010",
		b"11111010111011111110101011",
		b"11111010101011110010011010",
		b"11111010011011110111101100",
		b"11111010001100001110111111",
		b"11111001111100111000110010",
		b"11111001101101110101100000",
		b"11111001011111000101100100",
		b"11111001010000101001011010",
		b"11111001000010100001011100",
		b"11111000110100101110000011",
		b"11111000100111001111100111",
		b"11111000011010000110100000",
		b"11111000001101010011000100",
		b"11111000000000110101101010",
		b"11110111110100101110100110",
		b"11110111101000111110001011",
		b"11110111011101100100101111",
		b"11110111010010100010100001",
		b"11110111000111110111110101",
		b"11110110111101100100111010",
		b"11110110110011101010000001",
		b"11110110101010000111010111",
		b"11110110100000111101001010",
		b"11110110011000001011101000",
		b"11110110001111110010111100",
		b"11110110000111110011010001",
		b"11110110000000001100110010",
		b"11110101111000111111100111",
		b"11110101110010001011111001",
		b"11110101101011110001110000",
		b"11110101100101110001010001",
		b"11110101100000001010100010",
		b"11110101011010111101100111",
		b"11110101010110001010100101",
		b"11110101010001110001011110",
		b"11110101001101110010010011",
		b"11110101001010001101000111",
		b"11110101000111000001111000",
		b"11110101000100010000100110",
		b"11110101000001111001010000",
		b"11110100111111111011110001",
		b"11110100111110011000001000",
		b"11110100111101001110001111",
		b"11110100111100011110000010",
		b"11110100111100000111011001",
		b"11110100111100001010001110",
		b"11110100111100100110011010",
		b"11110100111101011011110011",
		b"11110100111110101010001111",
		b"11110101000000010001100101",
		b"11110101000010010001101010",
		b"11110101000100101010010000",
		b"11110101000111011011001100",
		b"11110101001010100100010000",
		b"11110101001110000101001101",
		b"11110101010001111101110100",
		b"11110101010110001101110110",
		b"11110101011010110101000001",
		b"11110101011111110011000110",
		b"11110101100101000111110000",
		b"11110101101010110010101110",
		b"11110101110000110011101100",
		b"11110101110111001010010110",
		b"11110101111101110110011000",
		b"11110110000100110111011011",
		b"11110110001100001101001010",
		b"11110110010011110111001110",
		b"11110110011011110101001111",
		b"11110110100100000110110110",
		b"11110110101100101011101010",
		b"11110110110101100011010011",
		b"11110110111110101101010110",
		b"11110111001000001001011010",
		b"11110111010001110111000100",
		b"11110111011011110101111000",
		b"11110111100110000101011100",
		b"11110111110000100101010011",
		b"11110111111011010101000001",
		b"11111000000110010100001001",
		b"11111000010001100010001101",
		b"11111000011100111110110000",
		b"11111000101000101001010100",
		b"11111000110100100001011010",
		b"11111001000000100110100011",
		b"11111001001100111000010001",
		b"11111001011001010110000100",
		b"11111001100101111111011100",
		b"11111001110010110011111010",
		b"11111001111111110010111101",
		b"11111010001100111100000101",
		b"11111010011010001110110000",
		b"11111010100111101010100000",
		b"11111010110101001110110001",
		b"11111011000010111011000100",
		b"11111011010000101110110111",
		b"11111011011110101001101000",
		b"11111011101100101010110110",
		b"11111011111010110010000000",
		b"11111100001000111110100011",
		b"11111100010111001111111111",
		b"11111100100101100101110001",
		b"11111100110011111111011000",
		b"11111101000010011100010010",
		b"11111101010000111011111101",
		b"11111101011111011101111000",
		b"11111101101110000001100001",
		b"11111101111100100110010111",
		b"11111110001011001011111000",
		b"11111110011001110001100100",
		b"11111110101000010110111000",
		b"11111110110110111011010100",
		b"11111111000101011110011000",
		b"11111111010011111111100010",
		b"11111111100010011110010010",
		b"11111111110000111010001000",
		b"11111111111111010010100101",
		b"00000000001101100111001000",
		b"00000000011011110111010001",
		b"00000000101010000010100011",
		b"00000000111000001000011110",
		b"00000001000110001000100011",
		b"00000001010100000010010101",
		b"00000001100001110101010101",
		b"00000001101111100001000111",
		b"00000001111101000101001100",
		b"00000010001010100001001001",
		b"00000010010111110100100000",
		b"00000010100100111110110111",
		b"00000010110001111111110010",
		b"00000010111110110110110101",
		b"00000011001011100011100110",
		b"00000011011000000101101011",
		b"00000011100100011100101011",
		b"00000011110000101000001101",
		b"00000011111100100111110111",
		b"00000100001000011011010010",
		b"00000100010100000010000110",
		b"00000100011111011011111100",
		b"00000100101010101000011110",
		b"00000100110101100111010110",
		b"00000101000000011000001111",
		b"00000101001010111010110011",
		b"00000101010101001110101111",
		b"00000101011111010011110000",
		b"00000101101001001001100001",
		b"00000101110010101111110001",
		b"00000101111100000110001111",
		b"00000110000101001100101000",
		b"00000110001110000010101101",
		b"00000110010110101000001110",
		b"00000110011110111100111011",
		b"00000110100111000000100110",
		b"00000110101110110011000010",
		b"00000110110110010100000000",
		b"00000110111101100011010101",
		b"00000111000100100000110100",
		b"00000111001011001100010011",
		b"00000111010001100101100111",
		b"00000111010111101100100101",
		b"00000111011101100001000110",
		b"00000111100011000011000000",
		b"00000111101000010010001011",
		b"00000111101101001110100010",
		b"00000111110001110111111100",
		b"00000111110110001110010101",
		b"00000111111010010001100111",
		b"00000111111110000001101110",
		b"00001000000001011110100111",
		b"00001000000100101000001110",
		b"00001000000111011110100010",
		b"00001000001010000001100000",
		b"00001000001100010001001000",
		b"00001000001110001101011010",
		b"00001000001111110110010110",
		b"00001000010001001011111101",
		b"00001000010010001110010010",
		b"00001000010010111101010110",
		b"00001000010011011001001110",
		b"00001000010011100001111011",
		b"00001000010011010111100101",
		b"00001000010010111010001110",
		b"00001000010010001001111110",
		b"00001000010001000110111011",
		b"00001000001111110001001011",
		b"00001000001110001000110111",
		b"00001000001100001110000111",
		b"00001000001010000001000100",
		b"00001000000111100001110111",
		b"00001000000100110000101010",
		b"00001000000001101101101001",
		b"00000111111110011000111111",
		b"00000111111010110010110111",
		b"00000111110110111011011111",
		b"00000111110010110011000011",
		b"00000111101110011001110000",
		b"00000111101001101111110110",
		b"00000111100100110101100010",
		b"00000111011111101011000100",
		b"00000111011010010000101100",
		b"00000111010100100110101010",
		b"00000111001110101101001110",
		b"00000111001000100100101010",
		b"00000111000010001101010000",
		b"00000110111011100111010001",
		b"00000110110100110011000000",
		b"00000110101101110000110000",
		b"00000110100110100000110101",
		b"00000110011111000011100010",
		b"00000110010111011001001100",
		b"00000110001111100010000111",
		b"00000110000111011110101000",
		b"00000101111111001111000101",
		b"00000101110110110011110011",
		b"00000101101110001101001000",
		b"00000101100101011011011010",
		b"00000101011100011111000001",
		b"00000101010011011000010011",
		b"00000101001010000111100111",
		b"00000101000000101101010101",
		b"00000100110111001001110101",
		b"00000100101101011101011110",
		b"00000100100011101000101001",
		b"00000100011001101011101110",
		b"00000100001111100111000110",
		b"00000100000101011011001001",
		b"00000011111011001000010000",
		b"00000011110000101110110101",
		b"00000011100110001111010001",
		b"00000011011011101001111101",
		b"00000011010000111111010010",
		b"00000011000110001111101010",
		b"00000010111011011011011111",
		b"00000010110000100011001011",
		b"00000010100101100111000111",
		b"00000010011010100111101100",
		b"00000010001111100101010110",
		b"00000010000100100000011101",
		b"00000001111001011001011011",
		b"00000001101110010000101011",
		b"00000001100011000110100110",
		b"00000001010111111011100101",
		b"00000001001100110000000011",
		b"00000001000001100100011001",
		b"00000000110110011001000000",
		b"00000000101011001110010010",
		b"00000000100000000100101000",
		b"00000000010100111100011100",
		b"00000000001001110110000101",
		b"11111111111110110001111110",
		b"11111111110011110000011110",
		b"11111111101000110001111111",
		b"11111111011101110110111001",
		b"11111111010010111111100011",
		b"11111111001000001100010101",
		b"11111110111101011101101000",
		b"11111110110010110011110010",
		b"11111110101000001111001100",
		b"11111110011101110000001010",
		b"11111110010011010111000101",
		b"11111110001001000100010010",
		b"11111101111110111000001000",
		b"11111101110100110010111100",
		b"11111101101010110101000011",
		b"11111101100000111110110011",
		b"11111101010111010000100001",
		b"11111101001101101010011111",
		b"11111101000100001101000011",
		b"11111100111010111000100001",
		b"11111100110001101101001010",
		b"11111100101000101011010011",
		b"11111100011111110011001101",
		b"11111100010111000101001010",
		b"11111100001110100001011101",
		b"11111100000110001000010110",
		b"11111011111101111010000101",
		b"11111011110101110110111100",
		b"11111011101101111111001010",
		b"11111011100110010010111110",
		b"11111011011110110010100111",
		b"11111011010111011110010100",
		b"11111011010000010110010010",
		b"11111011001001011010101111",
		b"11111011000010101011111001",
		b"11111010111100001001111010",
		b"11111010110101110101000001",
		b"11111010101111101101010111",
		b"11111010101001110011001000",
		b"11111010100100000110011110",
		b"11111010011110100111100011",
		b"11111010011001010110100001",
		b"11111010010100010011100001",
		b"11111010001111011110101010",
		b"11111010001010111000000101",
		b"11111010000110011111111001",
		b"11111010000010010110001101",
		b"11111001111110011011000111",
		b"11111001111010101110101100",
		b"11111001110111010001000010",
		b"11111001110100000010001101",
		b"11111001110001000010010010",
		b"11111001101110010001010100",
		b"11111001101011101111010110",
		b"11111001101001011100011010",
		b"11111001100111011000100010",
		b"11111001100101100011110000",
		b"11111001100011111110000100",
		b"11111001100010100111011111",
		b"11111001100001100000000000",
		b"11111001100000100111100111",
		b"11111001011111111110010010",
		b"11111001011111100011111111",
		b"11111001011111011000101101",
		b"11111001011111011100010111",
		b"11111001011111101110111011",
		b"11111001100000010000010101",
		b"11111001100001000000100001",
		b"11111001100001111111011000",
		b"11111001100011001100110111",
		b"11111001100100101000110110",
		b"11111001100110010011001111",
		b"11111001101000001011111100",
		b"11111001101010010010110110",
		b"11111001101100100111110011",
		b"11111001101111001010101100",
		b"11111001110001111011011000",
		b"11111001110100111001101101",
		b"11111001111000000101100010",
		b"11111001111011011110101101",
		b"11111001111111000101000010",
		b"11111010000010111000011000",
		b"11111010000110111000100010",
		b"11111010001011000101010100",
		b"11111010001111011110100011",
		b"11111010010100000100000001",
		b"11111010011000110101100001",
		b"11111010011101110010110110",
		b"11111010100010111011110010",
		b"11111010101000010000000111",
		b"11111010101101101111100110",
		b"11111010110011011010000000",
		b"11111010111001001111000101",
		b"11111010111111001110101000",
		b"11111011000101011000010110",
		b"11111011001011101100000001",
		b"11111011010010001001010111",
		b"11111011011000110000001000",
		b"11111011011111100000000011",
		b"11111011100110011000110110",
		b"11111011101101011010010000",
		b"11111011110100100011111110",
		b"11111011111011110101110000",
		b"11111100000011001111010010",
		b"11111100001010110000010010",
		b"11111100010010011000011101",
		b"11111100011010000111100000",
		b"11111100100001111101001000",
		b"11111100101001111001000010",
		b"11111100110001111010111011",
		b"11111100111010000010011110",
		b"11111101000010001111011000",
		b"11111101001010100001010110",
		b"11111101010010111000000011",
		b"11111101011011010011001011",
		b"11111101100011110010011010",
		b"11111101101100010101011100",
		b"11111101110100111011111100",
		b"11111101111101100101100111",
		b"11111110000110010010000111",
		b"11111110001111000001001000",
		b"11111110010111110010010111",
		b"11111110100000100101011101",
		b"11111110101001011010001000",
		b"11111110110010010000000010",
		b"11111110111011000110110111",
		b"11111111000011111110010010",
		b"11111111001100110110000000",
		b"11111111010101101101101100",
		b"11111111011110100101000001",
		b"11111111100111011011101100",
		b"11111111110000010001011000",
		b"11111111111001000101110010",
		b"00000000000001111000100110",
		b"00000000001010101001011111",
		b"00000000010011011000001011",
		b"00000000011100000100010110",
		b"00000000100100101101101100",
		b"00000000101101010011111011",
		b"00000000110101110110101111",
		b"00000000111110010101110110",
		b"00000001000110110000111101",
		b"00000001001111000111110001",
		b"00000001010111011010000010",
		b"00000001011111100111011100",
		b"00000001100111101111101101",
		b"00000001101111110010100101",
		b"00000001110111101111110010",
		b"00000001111111100111000100",
		b"00000010000111011000001000",
		b"00000010001111000010110000",
		b"00000010010110100110101011",
		b"00000010011110000011101001",
		b"00000010100101011001011010",
		b"00000010101100100111101111",
		b"00000010110011101110011001",
		b"00000010111010101101001011",
		b"00000011000001100011110100",
		b"00000011001000010010001000",
		b"00000011001110110111111000",
		b"00000011010101010100111000",
		b"00000011011011101000111010",
		b"00000011100001110011110011",
		b"00000011100111110101010101",
		b"00000011101101101101010101",
		b"00000011110011011011100111",
		b"00000011111001000000000001",
		b"00000011111110011010010111",
		b"00000100000011101010100001",
		b"00000100001000110000010010",
		b"00000100001101101011100011",
		b"00000100010010011100001010",
		b"00000100010111000001111110",
		b"00000100011011011100110111",
		b"00000100011111101100101101",
		b"00000100100011110001011001",
		b"00000100100111101010110011",
		b"00000100101011011000110110",
		b"00000100101110111011011011",
		b"00000100110010010010011100",
		b"00000100110101011101110011",
		b"00000100111000011101011101",
		b"00000100111011010001010101",
		b"00000100111101111001010110",
		b"00000101000000010101011101",
		b"00000101000010100101100111",
		b"00000101000100101001110001",
		b"00000101000110100001111000",
		b"00000101001000001101111100",
		b"00000101001001101101111011",
		b"00000101001011000001110011",
		b"00000101001100001001100100",
		b"00000101001101000101001110",
		b"00000101001101110100110010",
		b"00000101001110011000001111",
		b"00000101001110101111101000",
		b"00000101001110111010111101",
		b"00000101001110111010010010",
		b"00000101001110101101101000",
		b"00000101001110010101000010",
		b"00000101001101110000100011",
		b"00000101001101000000010000",
		b"00000101001100000100001100",
		b"00000101001010111100011100",
		b"00000101001001101001000100",
		b"00000101001000001010001011",
		b"00000101000110011111110101",
		b"00000101000100101010001001",
		b"00000101000010101001001101",
		b"00000101000000011101001000",
		b"00000100111110000110000010",
		b"00000100111011100100000010",
		b"00000100111000110111001111",
		b"00000100110101111111110011",
		b"00000100110010111101110110",
		b"00000100101111110001100001",
		b"00000100101100011010111101",
		b"00000100101000111010010100",
		b"00000100100101001111110001",
		b"00000100100001011011011100",
		b"00000100011101011101100010",
		b"00000100011001010110001100",
		b"00000100010101000101100111",
		b"00000100010000101011111110",
		b"00000100001100001001011101",
		b"00000100000111011110001111",
		b"00000100000010101010100010",
		b"00000011111101101110100010",
		b"00000011111000101010011011",
		b"00000011110011011110011011",
		b"00000011101110001010110000",
		b"00000011101000101111100111",
		b"00000011100011001101001110",
		b"00000011011101100011110011",
		b"00000011010111110011100100",
		b"00000011010001111100110000",
		b"00000011001011111111100101",
		b"00000011000101111100010011",
		b"00000010111111110011001000",
		b"00000010111001100100010100",
		b"00000010110011010000000101",
		b"00000010101100110110101100",
		b"00000010100110011000011000",
		b"00000010011111110101011000",
		b"00000010011001001101111101",
		b"00000010010010100010010111",
		b"00000010001011110010110101",
		b"00000010000100111111101000",
		b"00000001111110001001000000",
		b"00000001110111001111001110",
		b"00000001110000010010100001",
		b"00000001101001010011001011",
		b"00000001100010010001011011",
		b"00000001011011001101100011",
		b"00000001010100000111110010",
		b"00000001001101000000011001",
		b"00000001000101110111101010",
		b"00000000111110101101110011",
		b"00000000110111100011000111",
		b"00000000110000010111110110",
		b"00000000101001001100001111",
		b"00000000100010000000100100",
		b"00000000011010110101000100",
		b"00000000010011101010000001",
		b"00000000001100011111101011",
		b"00000000000101010110010001",
		b"11111111111110001110000100",
		b"11111111110111000111010100",
		b"11111111110000000010010000",
		b"11111111101000111111001010",
		b"11111111100001111110010000",
		b"11111111011010111111110010",
		b"11111111010100000011111111",
		b"11111111001101001011000111",
		b"11111111000110010101011001",
		b"11111110111111100011000100",
		b"11111110111000110100010110",
		b"11111110110010001001011111",
		b"11111110101011100010101101",
		b"11111110100101000000001110",
		b"11111110011110100010010001",
		b"11111110011000001001000010",
		b"11111110010001110100110001",
		b"11111110001011100101101001",
		b"11111110000101011011111001",
		b"11111101111111010111101110",
		b"11111101111001011001010100",
		b"11111101110011100000111000",
		b"11111101101101101110100110",
		b"11111101101000000010101010",
		b"11111101100010011101010000",
		b"11111101011100111110100100",
		b"11111101010111100110110000",
		b"11111101010010010101111111",
		b"11111101001101001100011101",
		b"11111101001000001010010011",
		b"11111101000011001111101100",
		b"11111100111110011100110001",
		b"11111100111001110001101100",
		b"11111100110101001110100110",
		b"11111100110000110011101000",
		b"11111100101100100000111010",
		b"11111100101000010110100101",
		b"11111100100100010100110001",
		b"11111100100000011011100100",
		b"11111100011100101011000111",
		b"11111100011001000011100000",
		b"11111100010101100100110101",
		b"11111100010010001111001110",
		b"11111100001111000010101111",
		b"11111100001011111111011111",
		b"11111100001001000101100010",
		b"11111100000110010100111110",
		b"11111100000011101101110111",
		b"11111100000001010000010000",
		b"11111011111110111100001111",
		b"11111011111100110001110110",
		b"11111011111010110001001000",
		b"11111011111000111010001001",
		b"11111011110111001100111010",
		b"11111011110101101001011101",
		b"11111011110100001111110101",
		b"11111011110011000000000010",
		b"11111011110001111010000110",
		b"11111011110000111110000001",
		b"11111011110000001011110100",
		b"11111011101111100011011110",
		b"11111011101111000100111110",
		b"11111011101110110000010101",
		b"11111011101110100101100000",
		b"11111011101110100100011111",
		b"11111011101110101101010000",
		b"11111011101110111111110000",
		b"11111011101111011011111101",
		b"11111011110000000001110100",
		b"11111011110000110001010010",
		b"11111011110001101010010011",
		b"11111011110010101100110100",
		b"11111011110011111000110000",
		b"11111011110101001110000011",
		b"11111011110110101100101000",
		b"11111011111000010100011010",
		b"11111011111010000101010011",
		b"11111011111011111111001110",
		b"11111011111110000010000101",
		b"11111100000000001101110001",
		b"11111100000010100010001011",
		b"11111100000100111111001101",
		b"11111100000111100100101111",
		b"11111100001010010010101010",
		b"11111100001101001000110111",
		b"11111100010000000111001100",
		b"11111100010011001101100010",
		b"11111100010110011011110000",
		b"11111100011001110001101101",
		b"11111100011101001111010001",
		b"11111100100000110100010001",
		b"11111100100100100000100101",
		b"11111100101000010100000010",
		b"11111100101100001110011110",
		b"11111100110000001111101111",
		b"11111100110100010111101100",
		b"11111100111000100110001000",
		b"11111100111100111010111001",
		b"11111101000001010101110100",
		b"11111101000101110110101110",
		b"11111101001010011101011100",
		b"11111101001111001001110001",
		b"11111101010011111011100010",
		b"11111101011000110010100100",
		b"11111101011101101110101001",
		b"11111101100010101111100110",
		b"11111101100111110101001110",
		b"11111101101100111111010101",
		b"11111101110010001101101111",
		b"11111101110111100000001110",
		b"11111101111100110110100110",
		b"11111110000010010000101001",
		b"11111110000111101110001011",
		b"11111110001101001110111111",
		b"11111110010010110010110111",
		b"11111110011000011001100110",
		b"11111110011110000010111111",
		b"11111110100011101110110101",
		b"11111110101001011100111001",
		b"11111110101111001100111111",
		b"11111110110100111110111001",
		b"11111110111010110010011001",
		b"11111111000000100111010010",
		b"11111111000110011101010110",
		b"11111111001100010100011001",
		b"11111111010010001100001011",
		b"11111111011000000100100000",
		b"11111111011101111101001010",
		b"11111111100011110101111100",
		b"11111111101001101110101000",
		b"11111111101111100111000000",
		b"11111111110101011110111000",
		b"11111111111011010110000010",
		b"00000000000001001100010001",
		b"00000000000111000001011000",
		b"00000000001100110101001001",
		b"00000000010010100111010111",
		b"00000000011000010111110110",
		b"00000000011110000110011001",
		b"00000000100011110010110011",
		b"00000000101001011100111000",
		b"00000000101111000100011010",
		b"00000000110100101001001111",
		b"00000000111010001011001000",
		b"00000000111111101001111011",
		b"00000001000101000101011011",
		b"00000001001010011101011101",
		b"00000001001111110001110101",
		b"00000001010101000010011000",
		b"00000001011010001110111010",
		b"00000001011111010111010000",
		b"00000001100100011011001111",
		b"00000001101001011010101100",
		b"00000001101110010101011110",
		b"00000001110011001011011001",
		b"00000001110111111100010011",
		b"00000001111100101000000011",
		b"00000010000001001110011111",
		b"00000010000101101111011101",
		b"00000010001010001010110011",
		b"00000010001110100000011010",
		b"00000010010010110000000111",
		b"00000010010110111001110011",
		b"00000010011010111101010101",
		b"00000010011110111010100101",
		b"00000010100010110001011011",
		b"00000010100110100001110000",
		b"00000010101010001011011011",
		b"00000010101101101110010111",
		b"00000010110001001010011100",
		b"00000010110100011111100011",
		b"00000010110111101101100110",
		b"00000010111010110100100000",
		b"00000010111101110100001010",
		b"00000011000000101100011111",
		b"00000011000011011101011010",
		b"00000011000110000110110110",
		b"00000011001000101000101110",
		b"00000011001011000010111101",
		b"00000011001101010101100000",
		b"00000011001111100000010011",
		b"00000011010001100011010011",
		b"00000011010011011110011011",
		b"00000011010101010001101010",
		b"00000011010110111100111100",
		b"00000011011000100000001111",
		b"00000011011001111011100010",
		b"00000011011011001110110001",
		b"00000011011100011001111101",
		b"00000011011101011101000011",
		b"00000011011110011000000011",
		b"00000011011111001010111100",
		b"00000011011111110101101110",
		b"00000011100000011000011000",
		b"00000011100000110010111100",
		b"00000011100001000101011001",
		b"00000011100001001111110001",
		b"00000011100001010010000100",
		b"00000011100001001100010100",
		b"00000011100000111110100011",
		b"00000011100000101000110010",
		b"00000011100000001011000100",
		b"00000011011111100101011011",
		b"00000011011110110111111011",
		b"00000011011110000010100110",
		b"00000011011101000101011111",
		b"00000011011100000000101011",
		b"00000011011010110100001100",
		b"00000011011001100000001000",
		b"00000011011000000100100011",
		b"00000011010110100001100000",
		b"00000011010100110111000110",
		b"00000011010011000101011001",
		b"00000011010001001100011110",
		b"00000011001111001100011100",
		b"00000011001101000101011000",
		b"00000011001010110111011001",
		b"00000011001000100010100100",
		b"00000011000110000111000000",
		b"00000011000011100100110100",
		b"00000011000000111100000111",
		b"00000010111110001101000000",
		b"00000010111011010111100111",
		b"00000010111000011100000011",
		b"00000010110101011010011100",
		b"00000010110010010010111010",
		b"00000010101111000101100101",
		b"00000010101011110010100110",
		b"00000010101000011010000101",
		b"00000010100100111100001011",
		b"00000010100001011001000001",
		b"00000010011101110000101111",
		b"00000010011010000011100000",
		b"00000010010110010001011100",
		b"00000010010010011010101101",
		b"00000010001110011111011101",
		b"00000010001010011111110101",
		b"00000010000110011011111111",
		b"00000010000010010100000110",
		b"00000001111110001000010011",
		b"00000001111001111000110001",
		b"00000001110101100101101010",
		b"00000001110001001111001001",
		b"00000001101100110101011000",
		b"00000001101000011000100001",
		b"00000001100011111000110000",
		b"00000001011111010110001111",
		b"00000001011010110001001010",
		b"00000001010110001001101010",
		b"00000001010001011111111100",
		b"00000001001100110100001010",
		b"00000001001000000110011110",
		b"00000001000011010111000101",
		b"00000000111110100110001010",
		b"00000000111001110011110111",
		b"00000000110101000000010111",
		b"00000000110000001011110110",
		b"00000000101011010110100000",
		b"00000000100110100000011110",
		b"00000000100001101001111101",
		b"00000000011100110011001000",
		b"00000000010111111100001001",
		b"00000000010011000101001100",
		b"00000000001110001110011100",
		b"00000000001001011000000100",
		b"00000000000100100010001110",
		b"11111111111111101101000111",
		b"11111111111010111000111000",
		b"11111111110110000101101101",
		b"11111111110001010011110000",
		b"11111111101100100011001100",
		b"11111111100111110100001100",
		b"11111111100011000110111010",
		b"11111111011110011011100001",
		b"11111111011001110010001010",
		b"11111111010101001011000001",
		b"11111111010000100110001110",
		b"11111111001100000011111101",
		b"11111111000111100100011000",
		b"11111111000011000111100111",
		b"11111110111110101101110100",
		b"11111110111010010111001010",
		b"11111110110110000011110001",
		b"11111110110001110011110010",
		b"11111110101101100111011000",
		b"11111110101001011110101001",
		b"11111110100101011001110001",
		b"11111110100001011000110110",
		b"11111110011101011100000010",
		b"11111110011001100011011100",
		b"11111110010101101111001101",
		b"11111110010001111111011101",
		b"11111110001110010100010011",
		b"11111110001010101101110111",
		b"11111110000111001100010000",
		b"11111110000011101111100110",
		b"11111110000000011000000000",
		b"11111101111101000101100011",
		b"11111101111001111000011000",
		b"11111101110110110000100011",
		b"11111101110011101110001100",
		b"11111101110000110001011000",
		b"11111101101101111010001101",
		b"11111101101011001000110000",
		b"11111101101000011101000111",
		b"11111101100101110111010111",
		b"11111101100011010111100100",
		b"11111101100000111101110100",
		b"11111101011110101010001011",
		b"11111101011100011100101100",
		b"11111101011010010101011011",
		b"11111101011000010100011110",
		b"11111101010110011001110110",
		b"11111101010100100101100111",
		b"11111101010010110111110100",
		b"11111101010001010000100000",
		b"11111101001111101111101101",
		b"11111101001110010101011110",
		b"11111101001101000001110100",
		b"11111101001011110100110010",
		b"11111101001010101110011001",
		b"11111101001001101110101010",
		b"11111101001000110101100110",
		b"11111101001000000011001111",
		b"11111101000111010111100100",
		b"11111101000110110010100110",
		b"11111101000110010100010101",
		b"11111101000101111100110010",
		b"11111101000101101011111011",
		b"11111101000101100001110000",
		b"11111101000101011110010000",
		b"11111101000101100001011011",
		b"11111101000101101011001110",
		b"11111101000101111011101000",
		b"11111101000110010010101000",
		b"11111101000110110000001011",
		b"11111101000111010100010000",
		b"11111101000111111110110011",
		b"11111101001000101111110010",
		b"11111101001001100111001010",
		b"11111101001010100100111001",
		b"11111101001011101000111010",
		b"11111101001100110011001010",
		b"11111101001110000011100101",
		b"11111101001111011010001000",
		b"11111101010000110110101110",
		b"11111101010010011001010011",
		b"11111101010100000001110010",
		b"11111101010101110000000110",
		b"11111101010111100100001011",
		b"11111101011001011101111011",
		b"11111101011011011101010001",
		b"11111101011101100010000111",
		b"11111101011111101100010111",
		b"11111101100001111011111101",
		b"11111101100100010000110001",
		b"11111101100110101010101101",
		b"11111101101001001001101011",
		b"11111101101011101101100101",
		b"11111101101110010110010011",
		b"11111101110001000011101111",
		b"11111101110011110101110010",
		b"11111101110110101100010100",
		b"11111101111001100111001111",
		b"11111101111100100110011010",
		b"11111101111111101001101111",
		b"11111110000010110001000101",
		b"11111110000101111100010101",
		b"11111110001001001011010111",
		b"11111110001100011110000010",
		b"11111110001111110100001111",
		b"11111110010011001101110101",
		b"11111110010110101010101100",
		b"11111110011010001010101011",
		b"11111110011101101101101010",
		b"11111110100001010011100001",
		b"11111110100100111100000110",
		b"11111110101000100111010001",
		b"11111110101100010100111001",
		b"11111110110000000100110100",
		b"11111110110011110110111011",
		b"11111110110111101011000100",
		b"11111110111011100001000110",
		b"11111110111111011000111000",
		b"11111111000011010010010001",
		b"11111111000111001101000111",
		b"11111111001011001001010010",
		b"11111111001111000110101000",
		b"11111111010011000101000000",
		b"11111111010111000100010000",
		b"11111111011011000100010000",
		b"11111111011111000100110110",
		b"11111111100011000101111001",
		b"11111111100111000111010000",
		b"11111111101011001000110001",
		b"11111111101111001010010100",
		b"11111111110011001011101111",
		b"11111111110111001100111000",
		b"11111111111011001101101000",
		b"11111111111111001101110100",
		b"00000000000011001101010101",
		b"00000000000111001100000000",
		b"00000000001011001001101100",
		b"00000000001111000110010010",
		b"00000000010011000001101000",
		b"00000000010110111011100110",
		b"00000000011010110100000011",
		b"00000000011110101010110101",
		b"00000000100010011111110110",
		b"00000000100110010010111100",
		b"00000000101010000011111111",
		b"00000000101101110010110111",
		b"00000000110001011111011100",
		b"00000000110101001001100101",
		b"00000000111000110001001011",
		b"00000000111100010110000111",
		b"00000000111111111000010000",
		b"00000001000011010111011110",
		b"00000001000110110011101011",
		b"00000001001010001100101111",
		b"00000001001101100010100100",
		b"00000001010000110101000001",
		b"00000001010100000100000000",
		b"00000001010111001111011011",
		b"00000001011010010111001010",
		b"00000001011101011011000111",
		b"00000001100000011011001101",
		b"00000001100011010111010100",
		b"00000001100110001111010111",
		b"00000001101001000011010001",
		b"00000001101011110010111010",
		b"00000001101110011110001111",
		b"00000001110001000101001001",
		b"00000001110011100111100100",
		b"00000001110110000101011010",
		b"00000001111000011110100111",
		b"00000001111010110011000101",
		b"00000001111101000010110010",
		b"00000001111111001101101000",
		b"00000010000001010011100011",
		b"00000010000011010100011111",
		b"00000010000101010000011010",
		b"00000010000111000111001110",
		b"00000010001000111000111010",
		b"00000010001010100101011001",
		b"00000010001100001100101001",
		b"00000010001101101110100111",
		b"00000010001111001011010001",
		b"00000010010000100010100100",
		b"00000010010001110100011111",
		b"00000010010011000000111110",
		b"00000010010100001000000001",
		b"00000010010101001001100110",
		b"00000010010110000101101011",
		b"00000010010110111100010000",
		b"00000010010111101101010011",
		b"00000010011000011000110100",
		b"00000010011000111110110010",
		b"00000010011001011111001101",
		b"00000010011001111010000101",
		b"00000010011010001111011001",
		b"00000010011010011111001010",
		b"00000010011010101001011001",
		b"00000010011010101110000101",
		b"00000010011010101101010001",
		b"00000010011010100110111100",
		b"00000010011010011011001001",
		b"00000010011010001001111000",
		b"00000010011001110011001011",
		b"00000010011001010111000011",
		b"00000010011000110101100100",
		b"00000010011000001110101111",
		b"00000010010111100010100110",
		b"00000010010110110001001100",
		b"00000010010101111010100100",
		b"00000010010100111110110000",
		b"00000010010011111101110011",
		b"00000010010010110111110010",
		b"00000010010001101100101111",
		b"00000010010000011100101101",
		b"00000010001111000111110001",
		b"00000010001101101101111110",
		b"00000010001100001111011001",
		b"00000010001010101100000110",
		b"00000010001001000100001000",
		b"00000010000111010111100110",
		b"00000010000101100110100010",
		b"00000010000011110001000011",
		b"00000010000001110111001101",
		b"00000001111111111001000101",
		b"00000001111101110110110001",
		b"00000001111011110000010110",
		b"00000001111001100101111001",
		b"00000001110111010111100000",
		b"00000001110101000101010001",
		b"00000001110010101111010010",
		b"00000001110000010101101001",
		b"00000001101101111000011011",
		b"00000001101011010111110000",
		b"00000001101000110011101101",
		b"00000001100110001100011001",
		b"00000001100011100001111011",
		b"00000001100000110100011001",
		b"00000001011110000011111001",
		b"00000001011011010000100011",
		b"00000001011000011010011110",
		b"00000001010101100001110000",
		b"00000001010010100110100001",
		b"00000001001111101000110111",
		b"00000001001100101000111010",
		b"00000001001001100110110010",
		b"00000001000110100010100100",
		b"00000001000011011100011010",
		b"00000001000000010100011001",
		b"00000000111101001010101010",
		b"00000000111001111111010101",
		b"00000000110110110010011111",
		b"00000000110011100100010010",
		b"00000000110000010100110101",
		b"00000000101101000100001111",
		b"00000000101001110010101000",
		b"00000000100110100000000111",
		b"00000000100011001100110101",
		b"00000000011111111000111000",
		b"00000000011100100100011001",
		b"00000000011001001111100000",
		b"00000000010101111010010011",
		b"00000000010010100100111010",
		b"00000000001111001111011110",
		b"00000000001011111010000101",
		b"00000000001000100100111000",
		b"00000000000101001111111101",
		b"00000000000001111011011101",
		b"11111111111110100111011111",
		b"11111111111011010100001010",
		b"11111111111000000001100101",
		b"11111111110100101111111001",
		b"11111111110001011111001011",
		b"11111111101110001111100101",
		b"11111111101011000001001100",
		b"11111111100111110100001000",
		b"11111111100100101000011111",
		b"11111111100001011110011010",
		b"11111111011110010101111110",
		b"11111111011011001111010011",
		b"11111111011000001010100000",
		b"11111111010101000111101010",
		b"11111111010010000110111001",
		b"11111111001111001000010011",
		b"11111111001100001011111110",
		b"11111111001001010010000001",
		b"11111111000110011010100010",
		b"11111111000011100101100111",
		b"11111111000000110011010110",
		b"11111110111110000011110101",
		b"11111110111011010111001001",
		b"11111110111000101101011000",
		b"11111110110110000110101000",
		b"11111110110011100010111110",
		b"11111110110001000010100000",
		b"11111110101110100101010001",
		b"11111110101100001011011001",
		b"11111110101001110100111010",
		b"11111110100111100001111011",
		b"11111110100101010010011111",
		b"11111110100011000110101011",
		b"11111110100000111110100011",
		b"11111110011110111010001100",
		b"11111110011100111001101010",
		b"11111110011010111101000000",
		b"11111110011001000100010010",
		b"11111110010111001111100100",
		b"11111110010101011110111010",
		b"11111110010011110010010101",
		b"11111110010010001001111010",
		b"11111110010000100101101100",
		b"11111110001111000101101101",
		b"11111110001101101010000000",
		b"11111110001100010010100111",
		b"11111110001010111111100101",
		b"11111110001001110000111100",
		b"11111110001000100110101110",
		b"11111110000111100000111101",
		b"11111110000110011111101010",
		b"11111110000101100010110111",
		b"11111110000100101010100101",
		b"11111110000011110110110110",
		b"11111110000011000111101010",
		b"11111110000010011101000011",
		b"11111110000001110111000001",
		b"11111110000001010101100100",
		b"11111110000000111000101101",
		b"11111110000000100000011100",
		b"11111110000000001100110001",
		b"11111101111111111101101100",
		b"11111101111111110011001101",
		b"11111101111111101101010011",
		b"11111101111111101011111101",
		b"11111101111111101111001100",
		b"11111101111111110110111101",
		b"11111110000000000011010000",
		b"11111110000000010100000011",
		b"11111110000000101001010110",
		b"11111110000001000011000110",
		b"11111110000001100001010001",
		b"11111110000010000011110111",
		b"11111110000010101010110101",
		b"11111110000011010110001000",
		b"11111110000100000101101111",
		b"11111110000100111001100110",
		b"11111110000101110001101100",
		b"11111110000110101101111110",
		b"11111110000111101110011000",
		b"11111110001000110010110111",
		b"11111110001001111011011001",
		b"11111110001011000111111010",
		b"11111110001100011000010111",
		b"11111110001101101100101100",
		b"11111110001111000100110101",
		b"11111110010000100000101111",
		b"11111110010010000000010101",
		b"11111110010011100011100100",
		b"11111110010101001010010111",
		b"11111110010110110100101011",
		b"11111110011000100010011010",
		b"11111110011010010011100000",
		b"11111110011100000111111000",
		b"11111110011101111111011111",
		b"11111110011111111010001110",
		b"11111110100001111000000001",
		b"11111110100011111000110100",
		b"11111110100101111100100000",
		b"11111110101000000011000001",
		b"11111110101010001100010001",
		b"11111110101100011000001011",
		b"11111110101110100110101010",
		b"11111110110000110111100111",
		b"11111110110011001010111111",
		b"11111110110101100000101001",
		b"11111110110111111000100010",
		b"11111110111010010010100100",
		b"11111110111100101110100111",
		b"11111110111111001100100111",
		b"11111111000001101100011101",
		b"11111111000100001110000100",
		b"11111111000110110001010110",
		b"11111111001001010110001011",
		b"11111111001011111100011111",
		b"11111111001110100100001011",
		b"11111111010001001101001001",
		b"11111111010011110111010010",
		b"11111111010110100010100001",
		b"11111111011001001110101110",
		b"11111111011011111011110101",
		b"11111111011110101001101101",
		b"11111111100001011000010010",
		b"11111111100100000111011101",
		b"11111111100110110111001000",
		b"11111111101001100111001011",
		b"11111111101100010111100001",
		b"11111111101111001000000100",
		b"11111111110001111000101101",
		b"11111111110100101001010110",
		b"11111111110111011001111001",
		b"11111111111010001010001111",
		b"11111111111100111010010010",
		b"11111111111111101001111101",
		b"00000000000010011001001000",
		b"00000000000101000111101110",
		b"00000000000111110101101001",
		b"00000000001010100010110010",
		b"00000000001101001111000100",
		b"00000000001111111010011000",
		b"00000000010010100100101001",
		b"00000000010101001101110001",
		b"00000000010111110101101010",
		b"00000000011010011100001111",
		b"00000000011101000001011001",
		b"00000000011111100101000011",
		b"00000000100010000111001000",
		b"00000000100100100111100010",
		b"00000000100111000110001011",
		b"00000000101001100011000000",
		b"00000000101011111101111001",
		b"00000000101110010110110010",
		b"00000000110000101101100110",
		b"00000000110011000010010001",
		b"00000000110101010100101100",
		b"00000000110111100100110100",
		b"00000000111001110010100011",
		b"00000000111011111101110110",
		b"00000000111110000110100111",
		b"00000001000000001100110010",
		b"00000001000010010000010011",
		b"00000001000100010001000110",
		b"00000001000110001111000111",
		b"00000001001000001010010001",
		b"00000001001010000010100001",
		b"00000001001011110111110011",
		b"00000001001101101010000100",
		b"00000001001111011001010000",
		b"00000001010001000101010011",
		b"00000001010010101110001011",
		b"00000001010100010011110100",
		b"00000001010101110110001011",
		b"00000001010111010101001110",
		b"00000001011000110000111001",
		b"00000001011010001001001010",
		b"00000001011011011101111111",
		b"00000001011100101111010101",
		b"00000001011101111101001001",
		b"00000001011111000111011011",
		b"00000001100000001110000111",
		b"00000001100001010001001100",
		b"00000001100010010000101000",
		b"00000001100011001100011001",
		b"00000001100100000100011111",
		b"00000001100100111000111000",
		b"00000001100101101001100010",
		b"00000001100110010110011101",
		b"00000001100110111111101000",
		b"00000001100111100101000010",
		b"00000001101000000110101010",
		b"00000001101000100100011111",
		b"00000001101000111110100011",
		b"00000001101001010100110011",
		b"00000001101001100111010001",
		b"00000001101001110101111100",
		b"00000001101010000000110100",
		b"00000001101010000111111010",
		b"00000001101010001011001110",
		b"00000001101010001010110001",
		b"00000001101010000110100011",
		b"00000001101001111110100110",
		b"00000001101001110010111001",
		b"00000001101001100011011111",
		b"00000001101001010000011001",
		b"00000001101000111001101000",
		b"00000001101000011111001101",
		b"00000001101000000001001010",
		b"00000001100111011111100001",
		b"00000001100110111010010011",
		b"00000001100110010001100011",
		b"00000001100101100101010011",
		b"00000001100100110101100100",
		b"00000001100100000010011010",
		b"00000001100011001011110111",
		b"00000001100010010001111101",
		b"00000001100001010100101111",
		b"00000001100000010100001111",
		b"00000001011111010000100001",
		b"00000001011110001001101000",
		b"00000001011100111111100110",
		b"00000001011011110010011111",
		b"00000001011010100010010111",
		b"00000001011001001111010000",
		b"00000001010111111001001110",
		b"00000001010110100000010101",
		b"00000001010101000100101000",
		b"00000001010011100110001011",
		b"00000001010010000101000011",
		b"00000001010000100001010010",
		b"00000001001110111010111101",
		b"00000001001101010010001000",
		b"00000001001011100110111000",
		b"00000001001001111001010000",
		b"00000001001000001001010100",
		b"00000001000110010111001010",
		b"00000001000100100010110110",
		b"00000001000010101100011011",
		b"00000001000000110100000000",
		b"00000000111110111001101000",
		b"00000000111100111101011000",
		b"00000000111010111111010100",
		b"00000000111000111111100011",
		b"00000000110110111110001000",
		b"00000000110100111011001000",
		b"00000000110010110110101000",
		b"00000000110000110000101110",
		b"00000000101110101001011110",
		b"00000000101100100000111110",
		b"00000000101010010111010001",
		b"00000000101000001100011111",
		b"00000000100110000000101010",
		b"00000000100011110011111010",
		b"00000000100001100110010010",
		b"00000000011111010111111001",
		b"00000000011101001000110011",
		b"00000000011010111001000101",
		b"00000000011000101000110101",
		b"00000000010110011000001000",
		b"00000000010100000111000011",
		b"00000000010001110101101011",
		b"00000000001111100100000101",
		b"00000000001101010010011000",
		b"00000000001011000000100111",
		b"00000000001000101110111000",
		b"00000000000110011101010001",
		b"00000000000100001011110101",
		b"00000000000001111010101011",
		b"11111111111111101001111000",
		b"11111111111101011001100000",
		b"11111111111011001001101001",
		b"11111111111000111010011000",
		b"11111111110110101011110001",
		b"11111111110100011101111001",
		b"11111111110010010000110110",
		b"11111111110000000100101101",
		b"11111111101101111001100001",
		b"11111111101011101111011000",
		b"11111111101001100110010110",
		b"11111111100111011110100001",
		b"11111111100101010111111100",
		b"11111111100011010010101100",
		b"11111111100001001110110110",
		b"11111111011111001100011111",
		b"11111111011101001011101001",
		b"11111111011011001100011010",
		b"11111111011001001110110111",
		b"11111111010111010011000010",
		b"11111111010101011001000000",
		b"11111111010011100000110110",
		b"11111111010001101010100110",
		b"11111111001111110110010101",
		b"11111111001110000100000111",
		b"11111111001100010011111111",
		b"11111111001010100110000000",
		b"11111111001000111010001111",
		b"11111111000111010000101111",
		b"11111111000101101001100011",
		b"11111111000100000100101101",
		b"11111111000010100010010010",
		b"11111111000001000010010101",
		b"11111110111111100100111000",
		b"11111110111110001001111101",
		b"11111110111100110001101001",
		b"11111110111011011011111101",
		b"11111110111010001000111101",
		b"11111110111000111000101001",
		b"11111110110111101011000110",
		b"11111110110110100000010101",
		b"11111110110101011000010111",
		b"11111110110100010011010000",
		b"11111110110011010001000001",
		b"11111110110010010001101100",
		b"11111110110001010101010010",
		b"11111110110000011011110110",
		b"11111110101111100101011000",
		b"11111110101110110001111011",
		b"11111110101110000001011110",
		b"11111110101101010100000100",
		b"11111110101100101001101101",
		b"11111110101100000010011011",
		b"11111110101011011110001110",
		b"11111110101010111101000111",
		b"11111110101010011111000110",
		b"11111110101010000100001101",
		b"11111110101001101100011010",
		b"11111110101001010111101111",
		b"11111110101001000110001100",
		b"11111110101000110111110001",
		b"11111110101000101100011101",
		b"11111110101000100100010001",
		b"11111110101000011111001100",
		b"11111110101000011101001101",
		b"11111110101000011110010101",
		b"11111110101000100010100011",
		b"11111110101000101001110110",
		b"11111110101000110100001100",
		b"11111110101001000001100110",
		b"11111110101001010010000010",
		b"11111110101001100101011111",
		b"11111110101001111011111011",
		b"11111110101010010101010110",
		b"11111110101010110001101101",
		b"11111110101011010001000000",
		b"11111110101011110011001101",
		b"11111110101100011000010001",
		b"11111110101101000000001100",
		b"11111110101101101010111010",
		b"11111110101110011000011011",
		b"11111110101111001000101011",
		b"11111110101111111011101001",
		b"11111110110000110001010011",
		b"11111110110001101001100101",
		b"11111110110010100100011110",
		b"11111110110011100001111011",
		b"11111110110100100001111001",
		b"11111110110101100100010101",
		b"11111110110110101001001101",
		b"11111110110111110000011110",
		b"11111110111000111010000101",
		b"11111110111010000101111111",
		b"11111110111011010100001000",
		b"11111110111100100100011110",
		b"11111110111101110110111101",
		b"11111110111111001011100010",
		b"11111111000000100010001001",
		b"11111111000001111010101111",
		b"11111111000011010101010001",
		b"11111111000100110001101011",
		b"11111111000110001111111001",
		b"11111111000111101111111001",
		b"11111111001001010001100100",
		b"11111111001010110100111010",
		b"11111111001100011001110100",
		b"11111111001110000000010000",
		b"11111111001111101000001010",
		b"11111111010001010001011101",
		b"11111111010010111100000110",
		b"11111111010100101000000001",
		b"11111111010110010101001001",
		b"11111111011000000011011011",
		b"11111111011001110010110010",
		b"11111111011011100011001010",
		b"11111111011101010100100000",
		b"11111111011111000110101110",
		b"11111111100000111001110001",
		b"11111111100010101101100101",
		b"11111111100100100010000101",
		b"11111111100110010111001101",
		b"11111111101000001100111000",
		b"11111111101010000011000011",
		b"11111111101011111001101010",
		b"11111111101101110000100111",
		b"11111111101111100111110111",
		b"11111111110001011111010101",
		b"11111111110011010110111110",
		b"11111111110101001110101100",
		b"11111111110111000110011100",
		b"11111111111000111110001001",
		b"11111111111010110101110000",
		b"11111111111100101101001100",
		b"11111111111110100100011000",
		b"00000000000000011011010001",
		b"00000000000010010001110011",
		b"00000000000100000111111001",
		b"00000000000101111101011111",
		b"00000000000111110010100010",
		b"00000000001001100110111100",
		b"00000000001011011010101011",
		b"00000000001101001101101011",
		b"00000000001110111111110110",
		b"00000000010000110001001011",
		b"00000000010010100001100011",
		b"00000000010100010000111101",
		b"00000000010101111111010100",
		b"00000000010111101100100100",
		b"00000000011001011000101010",
		b"00000000011011000011100011",
		b"00000000011100101101001001",
		b"00000000011110010101011011",
		b"00000000011111111100010101",
		b"00000000100001100001110011",
		b"00000000100011000101110011",
		b"00000000100100101000010000",
		b"00000000100110001001000111",
		b"00000000100111101000010111",
		b"00000000101001000101111010",
		b"00000000101010100001110000",
		b"00000000101011111011110011",
		b"00000000101101010100000011",
		b"00000000101110101010011011",
		b"00000000101111111110111010",
		b"00000000110001010001011101",
		b"00000000110010100010000001",
		b"00000000110011110000100011",
		b"00000000110100111101000010",
		b"00000000110110000111011010",
		b"00000000110111001111101011",
		b"00000000111000010101110001",
		b"00000000111001011001101011",
		b"00000000111010011011010110",
		b"00000000111011011010110001",
		b"00000000111100010111111010",
		b"00000000111101010010101111",
		b"00000000111110001011001111",
		b"00000000111111000001010111",
		b"00000000111111110101001000",
		b"00000001000000100110011110",
		b"00000001000001010101011010",
		b"00000001000010000001111001",
		b"00000001000010101011111011",
		b"00000001000011010011011110",
		b"00000001000011111000100010",
		b"00000001000100011011000110",
		b"00000001000100111011001010",
		b"00000001000101011000101011",
		b"00000001000101110011101011",
		b"00000001000110001100001000",
		b"00000001000110100010000010",
		b"00000001000110110101011010",
		b"00000001000111000110001101",
		b"00000001000111010100011110",
		b"00000001000111100000001011",
		b"00000001000111101001010100",
		b"00000001000111101111111010",
		b"00000001000111110011111110",
		b"00000001000111110101011110",
		b"00000001000111110100011101",
		b"00000001000111110000111010",
		b"00000001000111101010110110",
		b"00000001000111100010010010",
		b"00000001000111010111001110",
		b"00000001000111001001101011",
		b"00000001000110111001101011",
		b"00000001000110100111001110",
		b"00000001000110010010010101",
		b"00000001000101111011000011",
		b"00000001000101100001010111",
		b"00000001000101000101010011",
		b"00000001000100100110111010",
		b"00000001000100000110001011",
		b"00000001000011100011001010",
		b"00000001000010111101110111",
		b"00000001000010010110010100",
		b"00000001000001101100100100",
		b"00000001000001000000101000",
		b"00000001000000010010100001",
		b"00000000111111100010010011",
		b"00000000111110101111111111",
		b"00000000111101111011101000",
		b"00000000111101000101001111",
		b"00000000111100001100110111",
		b"00000000111011010010100010",
		b"00000000111010010110010011",
		b"00000000111001011000001100",
		b"00000000111000011000010000",
		b"00000000110111010110100010",
		b"00000000110110010011000011",
		b"00000000110101001101111000",
		b"00000000110100000111000001",
		b"00000000110010111110100100",
		b"00000000110001110100100001",
		b"00000000110000101000111101",
		b"00000000101111011011111001",
		b"00000000101110001101011010",
		b"00000000101100111101100010",
		b"00000000101011101100010100",
		b"00000000101010011001110100",
		b"00000000101001000110000100",
		b"00000000100111110001001000",
		b"00000000100110011011000011",
		b"00000000100101000011111000",
		b"00000000100011101011101010",
		b"00000000100010010010011101",
		b"00000000100000111000010101",
		b"00000000011111011101010011",
		b"00000000011110000001011101",
		b"00000000011100100100110101",
		b"00000000011011000111011110",
		b"00000000011001101001011101",
		b"00000000011000001010110100",
		b"00000000010110101011100111",
		b"00000000010101001011111010",
		b"00000000010011101011101111",
		b"00000000010010001011001011",
		b"00000000010000101010010001",
		b"00000000001111001001000100",
		b"00000000001101100111101000",
		b"00000000001100000110000000",
		b"00000000001010100100010000",
		b"00000000001001000010011011",
		b"00000000000111100000100101",
		b"00000000000101111110110001",
		b"00000000000100011101000011",
		b"00000000000010111011011101",
		b"00000000000001011010000100",
		b"11111111111111111000111011",
		b"11111111111110011000000101",
		b"11111111111100110111100101",
		b"11111111111011010111100000",
		b"11111111111001110111110111",
		b"11111111111000011000101111",
		b"11111111110110111010001010",
		b"11111111110101011100001101",
		b"11111111110011111110111001",
		b"11111111110010100010010011",
		b"11111111110001000110011101",
		b"11111111101111101011011010",
		b"11111111101110010001001110",
		b"11111111101100110111111011",
		b"11111111101011011111100101",
		b"11111111101010001000001110",
		b"11111111101000110001111001",
		b"11111111100111011100101010",
		b"11111111100110001000100010",
		b"11111111100100110101100101",
		b"11111111100011100011110101",
		b"11111111100010010011010101",
		b"11111111100001000100000111",
		b"11111111011111110110001111",
		b"11111111011110101001101110",
		b"11111111011101011110100111",
		b"11111111011100010100111100",
		b"11111111011011001100110000",
		b"11111111011010000110000100",
		b"11111111011001000000111100",
		b"11111111010111111101011001",
		b"11111111010110111011011101",
		b"11111111010101111011001010",
		b"11111111010100111100100011",
		b"11111111010011111111101000",
		b"11111111010011000100011100",
		b"11111111010010001011000001",
		b"11111111010001010011011000",
		b"11111111010000011101100011",
		b"11111111001111101001100011",
		b"11111111001110110111011010",
		b"11111111001110000111001001",
		b"11111111001101011000110010",
		b"11111111001100101100010101",
		b"11111111001100000001110101",
		b"11111111001011011001010001",
		b"11111111001010110010101100",
		b"11111111001010001110000110",
		b"11111111001001101011100000",
		b"11111111001001001010111010",
		b"11111111001000101100010110",
		b"11111111001000001111110101",
		b"11111111000111110101010110",
		b"11111111000111011100111010",
		b"11111111000111000110100011",
		b"11111111000110110010001111",
		b"11111111000110100000000000",
		b"11111111000110001111110110",
		b"11111111000110000001110000",
		b"11111111000101110101101111",
		b"11111111000101101011110100",
		b"11111111000101100011111101",
		b"11111111000101011110001011",
		b"11111111000101011010011101",
		b"11111111000101011000110100",
		b"11111111000101011001001111",
		b"11111111000101011011101101",
		b"11111111000101100000001110",
		b"11111111000101100110110001",
		b"11111111000101101111010110",
		b"11111111000101111001111100",
		b"11111111000110000110100011",
		b"11111111000110010101001001",
		b"11111111000110100101101101",
		b"11111111000110111000001111",
		b"11111111000111001100101110",
		b"11111111000111100011001000",
		b"11111111000111111011011100",
		b"11111111001000010101101001",
		b"11111111001000110001101110",
		b"11111111001001001111101001",
		b"11111111001001101111011001",
		b"11111111001010010000111101",
		b"11111111001010110100010010",
		b"11111111001011011001011000",
		b"11111111001100000000001100",
		b"11111111001100101000101101",
		b"11111111001101010010111010",
		b"11111111001101111110101111",
		b"11111111001110101100001101",
		b"11111111001111011011001111",
		b"11111111010000001011110110",
		b"11111111010000111101111110",
		b"11111111010001110001100101",
		b"11111111010010100110101010",
		b"11111111010011011101001010",
		b"11111111010100010101000100",
		b"11111111010101001110010100",
		b"11111111010110001000111000",
		b"11111111010111000100101111",
		b"11111111011000000001110101",
		b"11111111011001000000001001",
		b"11111111011001111111101000",
		b"11111111011011000000010000",
		b"11111111011100000001111101",
		b"11111111011101000100101110",
		b"11111111011110001000100001",
		b"11111111011111001101010001",
		b"11111111100000010010111101",
		b"11111111100001011001100011",
		b"11111111100010100000111111",
		b"11111111100011101001001110",
		b"11111111100100110010001111",
		b"11111111100101111011111110",
		b"11111111100111000110011001",
		b"11111111101000010001011101",
		b"11111111101001011101000111",
		b"11111111101010101001010101",
		b"11111111101011110110000011",
		b"11111111101101000011001110",
		b"11111111101110010000110101",
		b"11111111101111011110110100",
		b"11111111110000101101001001",
		b"11111111110001111011110000",
		b"11111111110011001010100110",
		b"11111111110100011001101010",
		b"11111111110101101000111000",
		b"11111111110110111000001101",
		b"11111111111000000111100111",
		b"11111111111001010111000010",
		b"11111111111010100110011100",
		b"11111111111011110101110011",
		b"11111111111101000101000011",
		b"11111111111110010100001001",
		b"11111111111111100011000011",
		b"00000000000000110001101111",
		b"00000000000010000000001001",
		b"00000000000011001110001110",
		b"00000000000100011011111101",
		b"00000000000101101001010010",
		b"00000000000110110110001011",
		b"00000000001000000010100101",
		b"00000000001001001110011110",
		b"00000000001010011001110011",
		b"00000000001011100100100001",
		b"00000000001100101110100111",
		b"00000000001101111000000001",
		b"00000000001111000000101101",
		b"00000000010000001000101001",
		b"00000000010001001111110010",
		b"00000000010010010110000110",
		b"00000000010011011011100011",
		b"00000000010100100000000111",
		b"00000000010101100011101110",
		b"00000000010110100110011000",
		b"00000000010111101000000010",
		b"00000000011000101000101001",
		b"00000000011001101000001101",
		b"00000000011010100110101010",
		b"00000000011011100011111111",
		b"00000000011100100000001010",
		b"00000000011101011011001001",
		b"00000000011110010100111010",
		b"00000000011111001101011100",
		b"00000000100000000100101100",
		b"00000000100000111010101010",
		b"00000000100001101111010010",
		b"00000000100010100010100101",
		b"00000000100011010100100000",
		b"00000000100100000101000010",
		b"00000000100100110100001001",
		b"00000000100101100001110100",
		b"00000000100110001110000010",
		b"00000000100110111000110010",
		b"00000000100111100010000010",
		b"00000000101000001001110001",
		b"00000000101000101111111110",
		b"00000000101001010100101001",
		b"00000000101001110111101111",
		b"00000000101010011001010001",
		b"00000000101010111001001101",
		b"00000000101011010111100010",
		b"00000000101011110100010001",
		b"00000000101100001111010111",
		b"00000000101100101000110101",
		b"00000000101101000000101010",
		b"00000000101101010110110110",
		b"00000000101101101011011000",
		b"00000000101101111110001111",
		b"00000000101110001111011100",
		b"00000000101110011110111101",
		b"00000000101110101100110100",
		b"00000000101110111000111111",
		b"00000000101111000011100000",
		b"00000000101111001100010100",
		b"00000000101111010011011110",
		b"00000000101111011000111100",
		b"00000000101111011100101111",
		b"00000000101111011110110111",
		b"00000000101111011111010101",
		b"00000000101111011110001001",
		b"00000000101111011011010010",
		b"00000000101111010110110010",
		b"00000000101111010000101010",
		b"00000000101111001000111001",
		b"00000000101110111111100000",
		b"00000000101110110100100000",
		b"00000000101110100111111001",
		b"00000000101110011001101101",
		b"00000000101110001001111100",
		b"00000000101101111000101000",
		b"00000000101101100101110000",
		b"00000000101101010001010110",
		b"00000000101100111011011011",
		b"00000000101100100100000001",
		b"00000000101100001011000111",
		b"00000000101011110000110000",
		b"00000000101011010100111101",
		b"00000000101010110111101111",
		b"00000000101010011001000110",
		b"00000000101001111001000110",
		b"00000000101001010111101110",
		b"00000000101000110101000001",
		b"00000000101000010000111111",
		b"00000000100111101011101011",
		b"00000000100111000101000111",
		b"00000000100110011101010010",
		b"00000000100101110100010000",
		b"00000000100101001010000010",
		b"00000000100100011110101010",
		b"00000000100011110010001001",
		b"00000000100011000100100001",
		b"00000000100010010101110101",
		b"00000000100001100110000101",
		b"00000000100000110101010100",
		b"00000000100000000011100100",
		b"00000000011111010000110111",
		b"00000000011110011101001110",
		b"00000000011101101000101100",
		b"00000000011100110011010010",
		b"00000000011011111101000011",
		b"00000000011011000110000001",
		b"00000000011010001110001110",
		b"00000000011001010101101011",
		b"00000000011000011100011100",
		b"00000000010111100010100010",
		b"00000000010110101000000000",
		b"00000000010101101100110110",
		b"00000000010100110001001001",
		b"00000000010011110100111010",
		b"00000000010010111000001011",
		b"00000000010001111010111110",
		b"00000000010000111101010110",
		b"00000000001111111111010101",
		b"00000000001111000000111101",
		b"00000000001110000010010000",
		b"00000000001101000011010001",
		b"00000000001100000100000010",
		b"00000000001011000100100100",
		b"00000000001010000100111100",
		b"00000000001001000101001010",
		b"00000000001000000101010001",
		b"00000000000111000101010011",
		b"00000000000110000101010010",
		b"00000000000101000101010010",
		b"00000000000100000101010011",
		b"00000000000011000101011000",
		b"00000000000010000101100011",
		b"00000000000001000101111000",
		b"00000000000000000110010110",
		b"11111111111111000111000010",
		b"11111111111110000111111101",
		b"11111111111101001001001001",
		b"11111111111100001010101001",
		b"11111111111011001100011110",
		b"11111111111010001110101010",
		b"11111111111001010001010001",
		b"11111111111000010100010011",
		b"11111111110111010111110010",
		b"11111111110110011011110010",
		b"11111111110101100000010011",
		b"11111111110100100101011000",
		b"11111111110011101011000011",
		b"11111111110010110001010101",
		b"11111111110001111000010001",
		b"11111111110000111111111000",
		b"11111111110000001000001100",
		b"11111111101111010001001111",
		b"11111111101110011011000011",
		b"11111111101101100101101001",
		b"11111111101100110001000100",
		b"11111111101011111101010100",
		b"11111111101011001010011011",
		b"11111111101010011000011100",
		b"11111111101001100111010111",
		b"11111111101000110111001110",
		b"11111111101000001000000011",
		b"11111111100111011001110110",
		b"11111111100110101100101010",
		b"11111111100110000000100000",
		b"11111111100101010101011001",
		b"11111111100100101011010110",
		b"11111111100100000010011001",
		b"11111111100011011010100010",
		b"11111111100010110011110100",
		b"11111111100010001110001110",
		b"11111111100001101001110011",
		b"11111111100001000110100011",
		b"11111111100000100100011111",
		b"11111111100000000011101000",
		b"11111111011111100011111111",
		b"11111111011111000101100100",
		b"11111111011110101000011010",
		b"11111111011110001100011111",
		b"11111111011101110001110110",
		b"11111111011101011000011111",
		b"11111111011101000000011001",
		b"11111111011100101001100111",
		b"11111111011100010100001000",
		b"11111111011011111111111101",
		b"11111111011011101101000110",
		b"11111111011011011011100100",
		b"11111111011011001011010111",
		b"11111111011010111100011111",
		b"11111111011010101110111100",
		b"11111111011010100010110000",
		b"11111111011010010111111001",
		b"11111111011010001110011000",
		b"11111111011010000110001101",
		b"11111111011001111111011000",
		b"11111111011001111001111001",
		b"11111111011001110101110000",
		b"11111111011001110010111100",
		b"11111111011001110001011110",
		b"11111111011001110001010110",
		b"11111111011001110010100010",
		b"11111111011001110101000011",
		b"11111111011001111000111000",
		b"11111111011001111110000001",
		b"11111111011010000100011110",
		b"11111111011010001100001101",
		b"11111111011010010101001111",
		b"11111111011010011111100011",
		b"11111111011010101011000111",
		b"11111111011010110111111101",
		b"11111111011011000110000010",
		b"11111111011011010101010110",
		b"11111111011011100101111000",
		b"11111111011011110111100111",
		b"11111111011100001010100011",
		b"11111111011100011110101011",
		b"11111111011100110011111101",
		b"11111111011101001010011001",
		b"11111111011101100001111110",
		b"11111111011101111010101010",
		b"11111111011110010100011100",
		b"11111111011110101111010100",
		b"11111111011111001011010000",
		b"11111111011111101000001111",
		b"11111111100000000110001111",
		b"11111111100000100101010000",
		b"11111111100001000101010000",
		b"11111111100001100110001110",
		b"11111111100010001000001001",
		b"11111111100010101010111110",
		b"11111111100011001110101101",
		b"11111111100011110011010101",
		b"11111111100100011000110011",
		b"11111111100100111111000111",
		b"11111111100101100110001110",
		b"11111111100110001110001000",
		b"11111111100110110110110010",
		b"11111111100111100000001011",
		b"11111111101000001010010010",
		b"11111111101000110101000101",
		b"11111111101001100000100010",
		b"11111111101010001100101000",
		b"11111111101010111001010100",
		b"11111111101011100110100110",
		b"11111111101100010100011100",
		b"11111111101101000010110011",
		b"11111111101101110001101010",
		b"11111111101110100001000000",
		b"11111111101111010000110010",
		b"11111111110000000001000000",
		b"11111111110000110001100110",
		b"11111111110001100010100100",
		b"11111111110010010011110111",
		b"11111111110011000101011110",
		b"11111111110011110111010111",
		b"11111111110100101001100001",
		b"11111111110101011011111000",
		b"11111111110110001110011101",
		b"11111111110111000001001100",
		b"11111111110111110100000100",
		b"11111111111000100111000011",
		b"11111111111001011010001000",
		b"11111111111010001101010000",
		b"11111111111011000000011010",
		b"11111111111011110011100101",
		b"11111111111100100110101101",
		b"11111111111101011001110010",
		b"11111111111110001100110010",
		b"11111111111110111111101010",
		b"11111111111111110010011010",
		b"00000000000000100101000000",
		b"00000000000001010111011001",
		b"00000000000010001001100100",
		b"00000000000010111011100000",
		b"00000000000011101101001010",
		b"00000000000100011110100010",
		b"00000000000101001111100101",
		b"00000000000110000000010010",
		b"00000000000110110000100110",
		b"00000000000111100000100010",
		b"00000000001000010000000010",
		b"00000000001000111111000110",
		b"00000000001001101101101011",
		b"00000000001010011011110001",
		b"00000000001011001001010110",
		b"00000000001011110110011001",
		b"00000000001100100010110111",
		b"00000000001101001110110000",
		b"00000000001101111010000010",
		b"00000000001110100100101100",
		b"00000000001111001110101100",
		b"00000000001111111000000001",
		b"00000000010000100000101010",
		b"00000000010001001000100110",
		b"00000000010001101111110011",
		b"00000000010010010110010001",
		b"00000000010010111011111101",
		b"00000000010011100000110111",
		b"00000000010100000100111110",
		b"00000000010100101000010001",
		b"00000000010101001010101110",
		b"00000000010101101100010100",
		b"00000000010110001101000100",
		b"00000000010110101100111011",
		b"00000000010111001011111001",
		b"00000000010111101001111100",
		b"00000000011000000111000101",
		b"00000000011000100011010010",
		b"00000000011000111110100011",
		b"00000000011001011000110110",
		b"00000000011001110010001011",
		b"00000000011010001010100001",
		b"00000000011010100001111001",
		b"00000000011010111000010000",
		b"00000000011011001101100111",
		b"00000000011011100001111101",
		b"00000000011011110101010010",
		b"00000000011100000111100101",
		b"00000000011100011000110101",
		b"00000000011100101001000011",
		b"00000000011100111000001110",
		b"00000000011101000110010110",
		b"00000000011101010011011010",
		b"00000000011101011111011010",
		b"00000000011101101010010111",
		b"00000000011101110100001111",
		b"00000000011101111101000011",
		b"00000000011110000100110011",
		b"00000000011110001011011111",
		b"00000000011110010001000110",
		b"00000000011110010101101001",
		b"00000000011110011001001000",
		b"00000000011110011011100011",
		b"00000000011110011100111010",
		b"00000000011110011101001101",
		b"00000000011110011100011101",
		b"00000000011110011010101001",
		b"00000000011110010111110011",
		b"00000000011110010011111010",
		b"00000000011110001110111111",
		b"00000000011110001001000010",
		b"00000000011110000010000011",
		b"00000000011101111010000011",
		b"00000000011101110001000011",
		b"00000000011101100111000100",
		b"00000000011101011100000100",
		b"00000000011101010000000110",
		b"00000000011101000011001010",
		b"00000000011100110101010001",
		b"00000000011100100110011010",
		b"00000000011100010110101000",
		b"00000000011100000101111010",
		b"00000000011011110100010010",
		b"00000000011011100001110000",
		b"00000000011011001110010101",
		b"00000000011010111010000010",
		b"00000000011010100100111001",
		b"00000000011010001110111000",
		b"00000000011001111000000011",
		b"00000000011001100000011010",
		b"00000000011001000111111101",
		b"00000000011000101110101110",
		b"00000000011000010100101110",
		b"00000000010111111001111101",
		b"00000000010111011110011110",
		b"00000000010111000010010001",
		b"00000000010110100101010111",
		b"00000000010110000111110001",
		b"00000000010101101001100001",
		b"00000000010101001010101000",
		b"00000000010100101011000110",
		b"00000000010100001010111110",
		b"00000000010011101010010000",
		b"00000000010011001000111110",
		b"00000000010010100111001000",
		b"00000000010010000100110001",
		b"00000000010001100001111010",
		b"00000000010000111110100011",
		b"00000000010000011010101111",
		b"00000000001111110110011110",
		b"00000000001111010001110010",
		b"00000000001110101100101100",
		b"00000000001110000111001110",
		b"00000000001101100001011001",
		b"00000000001100111011001110",
		b"00000000001100010100101111",
		b"00000000001011101101111110",
		b"00000000001011000110111010",
		b"00000000001010011111100111",
		b"00000000001001111000000101",
		b"00000000001001010000010110",
		b"00000000001000101000011011",
		b"00000000001000000000010110",
		b"00000000000111011000001000",
		b"00000000000110101111110010",
		b"00000000000110000111010110",
		b"00000000000101011110110110",
		b"00000000000100110110010010",
		b"00000000000100001101101100",
		b"00000000000011100101000110",
		b"00000000000010111100100001",
		b"00000000000010010011111110",
		b"00000000000001101011011111",
		b"00000000000001000011000101",
		b"00000000000000011010110001",
		b"11111111111111110010100101",
		b"11111111111111001010100011",
		b"11111111111110100010101011",
		b"11111111111101111010111111",
		b"11111111111101010011100000",
		b"11111111111100101100001111",
		b"11111111111100000101001111",
		b"11111111111011011110011111",
		b"11111111111010111000000010",
		b"11111111111010010001111001",
		b"11111111111001101100000101",
		b"11111111111001000110100110",
		b"11111111111000100001011111",
		b"11111111110111111100110001",
		b"11111111110111011000011100",
		b"11111111110110110100100010",
		b"11111111110110010001000100",
		b"11111111110101101110000011",
		b"11111111110101001011100001",
		b"11111111110100101001011101",
		b"11111111110100000111111011",
		b"11111111110011100110111001",
		b"11111111110011000110011010",
		b"11111111110010100110011111",
		b"11111111110010000111000111",
		b"11111111110001101000010110",
		b"11111111110001001010001010",
		b"11111111110000101100100110",
		b"11111111110000001111101010",
		b"11111111101111110011010110",
		b"11111111101111010111101101",
		b"11111111101110111100101110",
		b"11111111101110100010011010",
		b"11111111101110001000110011",
		b"11111111101101101111111000",
		b"11111111101101010111101011",
		b"11111111101101000000001100",
		b"11111111101100101001011011",
		b"11111111101100010011011011",
		b"11111111101011111110001010",
		b"11111111101011101001101010",
		b"11111111101011010101111011",
		b"11111111101011000010111101",
		b"11111111101010110000110010",
		b"11111111101010011111011001",
		b"11111111101010001110110100",
		b"11111111101001111111000001",
		b"11111111101001110000000010",
		b"11111111101001100001111000",
		b"11111111101001010100100010",
		b"11111111101001001000000000",
		b"11111111101000111100010011",
		b"11111111101000110001011011",
		b"11111111101000100111011001",
		b"11111111101000011110001100",
		b"11111111101000010101110100",
		b"11111111101000001110010011",
		b"11111111101000000111100110",
		b"11111111101000000001110000",
		b"11111111100111111100110000",
		b"11111111100111111000100101",
		b"11111111100111110101001111",
		b"11111111100111110010110000",
		b"11111111100111110001000110",
		b"11111111100111110000010001",
		b"11111111100111110000010010",
		b"11111111100111110001000111",
		b"11111111100111110010110010",
		b"11111111100111110101010001",
		b"11111111100111111000100100",
		b"11111111100111111100101011",
		b"11111111101000000001100110",
		b"11111111101000000111010100",
		b"11111111101000001101110101",
		b"11111111101000010101001001",
		b"11111111101000011101001111",
		b"11111111101000100110000110",
		b"11111111101000101111101110",
		b"11111111101000111010000111",
		b"11111111101001000101010001",
		b"11111111101001010001001001",
		b"11111111101001011101110001",
		b"11111111101001101011000111",
		b"11111111101001111001001011",
		b"11111111101010000111111100",
		b"11111111101010010111011010",
		b"11111111101010100111100011",
		b"11111111101010111000010111",
		b"11111111101011001001110101",
		b"11111111101011011011111101",
		b"11111111101011101110101110",
		b"11111111101100000010000111",
		b"11111111101100010110000111",
		b"11111111101100101010101101",
		b"11111111101100111111111001",
		b"11111111101101010101101010",
		b"11111111101101101011111110",
		b"11111111101110000010110101",
		b"11111111101110011010001110",
		b"11111111101110110010001000",
		b"11111111101111001010100010",
		b"11111111101111100011011100",
		b"11111111101111111100110011",
		b"11111111110000010110101000",
		b"11111111110000110000111001",
		b"11111111110001001011100101",
		b"11111111110001100110101100",
		b"11111111110010000010001011",
		b"11111111110010011110000011",
		b"11111111110010111010010010",
		b"11111111110011010110110110",
		b"11111111110011110011110000",
		b"11111111110100010000111110",
		b"11111111110100101110011111",
		b"11111111110101001100010001",
		b"11111111110101101010010100",
		b"11111111110110001000100110",
		b"11111111110110100111001000",
		b"11111111110111000101110110",
		b"11111111110111100100110001",
		b"11111111111000000011110111",
		b"11111111111000100011000111",
		b"11111111111001000010100000",
		b"11111111111001100010000001",
		b"11111111111010000001101000",
		b"11111111111010100001010110",
		b"11111111111011000001001000",
		b"11111111111011100000111101",
		b"11111111111100000000110101",
		b"11111111111100100000101101",
		b"11111111111101000000100110",
		b"11111111111101100000011110",
		b"11111111111110000000010100",
		b"11111111111110100000000111",
		b"11111111111110111111110110",
		b"11111111111111011111011111",
		b"11111111111111111111000010",
		b"00000000000000011110011110",
		b"00000000000000111101110001",
		b"00000000000001011100111011",
		b"00000000000001111011111010",
		b"00000000000010011010101110",
		b"00000000000010111001010101",
		b"00000000000011010111101111",
		b"00000000000011110101111010",
		b"00000000000100010011110101",
		b"00000000000100110001100000",
		b"00000000000101001110111010",
		b"00000000000101101100000001",
		b"00000000000110001000110100",
		b"00000000000110100101010100",
		b"00000000000111000001011110",
		b"00000000000111011101010011",
		b"00000000000111111000110000",
		b"00000000001000010011110110",
		b"00000000001000101110100011",
		b"00000000001001001000110110",
		b"00000000001001100010110000",
		b"00000000001001111100001110",
		b"00000000001010010101010000",
		b"00000000001010101101110110",
		b"00000000001011000101111111",
		b"00000000001011011101101010",
		b"00000000001011110100110110",
		b"00000000001100001011100010",
		b"00000000001100100001101111",
		b"00000000001100110111011010",
		b"00000000001101001100100101",
		b"00000000001101100001001101",
		b"00000000001101110101010011",
		b"00000000001110001000110110",
		b"00000000001110011011110101",
		b"00000000001110101110010000",
		b"00000000001111000000000110",
		b"00000000001111010001011000",
		b"00000000001111100010000011",
		b"00000000001111110010001001",
		b"00000000010000000001101000",
		b"00000000010000010000100001",
		b"00000000010000011110110010",
		b"00000000010000101100011100",
		b"00000000010000111001011110",
		b"00000000010001000101110111",
		b"00000000010001010001101001",
		b"00000000010001011100110001",
		b"00000000010001100111010001",
		b"00000000010001110001000111",
		b"00000000010001111010010100",
		b"00000000010010000010111000",
		b"00000000010010001010110010",
		b"00000000010010010010000010",
		b"00000000010010011000101001",
		b"00000000010010011110100101",
		b"00000000010010100011111000",
		b"00000000010010101000100000",
		b"00000000010010101100011110",
		b"00000000010010101111110011",
		b"00000000010010110010011101",
		b"00000000010010110100011110",
		b"00000000010010110101110101",
		b"00000000010010110110100010",
		b"00000000010010110110100101",
		b"00000000010010110101111111",
		b"00000000010010110100101111",
		b"00000000010010110010110111",
		b"00000000010010110000010110",
		b"00000000010010101101001100",
		b"00000000010010101001011001",
		b"00000000010010100100111111",
		b"00000000010010011111111100",
		b"00000000010010011010010011",
		b"00000000010010010100000001",
		b"00000000010010001101001010",
		b"00000000010010000101101011",
		b"00000000010001111101100111",
		b"00000000010001110100111101",
		b"00000000010001101011101110",
		b"00000000010001100001111001",
		b"00000000010001010111100001",
		b"00000000010001001100100101",
		b"00000000010001000001000101",
		b"00000000010000110101000011",
		b"00000000010000101000011110",
		b"00000000010000011011011000",
		b"00000000010000001101110000",
		b"00000000001111111111101000",
		b"00000000001111110001000000",
		b"00000000001111100001111001",
		b"00000000001111010010010011",
		b"00000000001111000010001110",
		b"00000000001110110001101100",
		b"00000000001110100000101110",
		b"00000000001110001111010011",
		b"00000000001101111101011101",
		b"00000000001101101011001100",
		b"00000000001101011000100001",
		b"00000000001101000101011101",
		b"00000000001100110010000001",
		b"00000000001100011110001100",
		b"00000000001100001010000001",
		b"00000000001011110101011111",
		b"00000000001011100000101000",
		b"00000000001011001011011100",
		b"00000000001010110101111100",
		b"00000000001010100000001001",
		b"00000000001010001010000100",
		b"00000000001001110011101101",
		b"00000000001001011101000101",
		b"00000000001001000110001110",
		b"00000000001000101111001000",
		b"00000000001000010111110011",
		b"00000000001000000000010001",
		b"00000000000111101000100011",
		b"00000000000111010000101001",
		b"00000000000110111000100100",
		b"00000000000110100000010110",
		b"00000000000110000111111110",
		b"00000000000101101111011110",
		b"00000000000101010110110110",
		b"00000000000100111110001000",
		b"00000000000100100101010100",
		b"00000000000100001100011100",
		b"00000000000011110011100000",
		b"00000000000011011010100000",
		b"00000000000011000001011110",
		b"00000000000010101000011011",
		b"00000000000010001111011000",
		b"00000000000001110110010100",
		b"00000000000001011101010010",
		b"00000000000001000100010010",
		b"00000000000000101011010101",
		b"00000000000000010010011011",
		b"11111111111111111001100110",
		b"11111111111111100000110110",
		b"11111111111111001000001100",
		b"11111111111110101111101010",
		b"11111111111110010111001111",
		b"11111111111101111110111100",
		b"11111111111101100110110011",
		b"11111111111101001110110100",
		b"11111111111100110111000000",
		b"11111111111100011111011000",
		b"11111111111100000111111100",
		b"11111111111011110000101101",
		b"11111111111011011001101100",
		b"11111111111011000010111001",
		b"11111111111010101100010110",
		b"11111111111010010110000011",
		b"11111111111010000000000001",
		b"11111111111001101010010000",
		b"11111111111001010100110001",
		b"11111111111000111111100101",
		b"11111111111000101010101100",
		b"11111111111000010110000111",
		b"11111111111000000001110111",
		b"11111111110111101101111100",
		b"11111111110111011010010111",
		b"11111111110111000111001000",
		b"11111111110110110100010000",
		b"11111111110110100001110000",
		b"11111111110110001111101000",
		b"11111111110101111101111000",
		b"11111111110101101100100001",
		b"11111111110101011011100100",
		b"11111111110101001011000001",
		b"11111111110100111010111001",
		b"11111111110100101011001011",
		b"11111111110100011011111001",
		b"11111111110100001101000011",
		b"11111111110011111110101001",
		b"11111111110011110000101011",
		b"11111111110011100011001011",
		b"11111111110011010110000111",
		b"11111111110011001001100010",
		b"11111111110010111101011010",
		b"11111111110010110001110000",
		b"11111111110010100110100101",
		b"11111111110010011011111001",
		b"11111111110010010001101011",
		b"11111111110010000111111101",
		b"11111111110001111110101111",
		b"11111111110001110110000000",
		b"11111111110001101101110000",
		b"11111111110001100110000001",
		b"11111111110001011110110010",
		b"11111111110001011000000011",
		b"11111111110001010001110101",
		b"11111111110001001100000111",
		b"11111111110001000110111001",
		b"11111111110001000010001100",
		b"11111111110000111110000000",
		b"11111111110000111010010100",
		b"11111111110000110111001001",
		b"11111111110000110100011110",
		b"11111111110000110010010100",
		b"11111111110000110000101011",
		b"11111111110000101111100010",
		b"11111111110000101110111001",
		b"11111111110000101110110000",
		b"11111111110000101111001000",
		b"11111111110000110000000000",
		b"11111111110000110001011000",
		b"11111111110000110011001111",
		b"11111111110000110101100110",
		b"11111111110000111000011100",
		b"11111111110000111011110001",
		b"11111111110000111111100101",
		b"11111111110001000011111000",
		b"11111111110001001000101010",
		b"11111111110001001101111001",
		b"11111111110001010011100110",
		b"11111111110001011001110001",
		b"11111111110001100000011000",
		b"11111111110001100111011101",
		b"11111111110001101110111110",
		b"11111111110001110110111100",
		b"11111111110001111111010101",
		b"11111111110010001000001010",
		b"11111111110010010001011001",
		b"11111111110010011011000011",
		b"11111111110010100101001000",
		b"11111111110010101111100110",
		b"11111111110010111010011101",
		b"11111111110011000101101101",
		b"11111111110011010001010110",
		b"11111111110011011101010110",
		b"11111111110011101001101110",
		b"11111111110011110110011100",
		b"11111111110100000011100001",
		b"11111111110100010000111100",
		b"11111111110100011110101100",
		b"11111111110100101100110001",
		b"11111111110100111011001010",
		b"11111111110101001001110110",
		b"11111111110101011000110110",
		b"11111111110101101000001000",
		b"11111111110101110111101101",
		b"11111111110110000111100010",
		b"11111111110110010111101000",
		b"11111111110110100111111110",
		b"11111111110110111000100100",
		b"11111111110111001001011001",
		b"11111111110111011010011100",
		b"11111111110111101011101101",
		b"11111111110111111101001010",
		b"11111111111000001110110100",
		b"11111111111000100000101010",
		b"11111111111000110010101011",
		b"11111111111001000100110110",
		b"11111111111001010111001011",
		b"11111111111001101001101010",
		b"11111111111001111100010000",
		b"11111111111010001110111111",
		b"11111111111010100001110101",
		b"11111111111010110100110001",
		b"11111111111011000111110011",
		b"11111111111011011010111010",
		b"11111111111011101110000110",
		b"11111111111100000001010110",
		b"11111111111100010100101001",
		b"11111111111100100111111110",
		b"11111111111100111011010101",
		b"11111111111101001110101110",
		b"11111111111101100010000111",
		b"11111111111101110101100000",
		b"11111111111110001000111000",
		b"11111111111110011100001111",
		b"11111111111110101111100100",
		b"11111111111111000010110110",
		b"11111111111111010110000101",
		b"11111111111111101001010000",
		b"11111111111111111100010110",
		b"00000000000000001111010111",
		b"00000000000000100010010010",
		b"00000000000000110101000111",
		b"00000000000001000111110101",
		b"00000000000001011010011011",
		b"00000000000001101100111000",
		b"00000000000001111111001101",
		b"00000000000010010001011001",
		b"00000000000010100011011010",
		b"00000000000010110101010001",
		b"00000000000011000110111101",
		b"00000000000011011000011101",
		b"00000000000011101001110000",
		b"00000000000011111010110111",
		b"00000000000100001011110001",
		b"00000000000100011100011100",
		b"00000000000100101100111010",
		b"00000000000100111101001000",
		b"00000000000101001101000111",
		b"00000000000101011100110111",
		b"00000000000101101100010110",
		b"00000000000101111011100100",
		b"00000000000110001010100001",
		b"00000000000110011001001100",
		b"00000000000110100111100101",
		b"00000000000110110101101100",
		b"00000000000111000011100000",
		b"00000000000111010001000000",
		b"00000000000111011110001101",
		b"00000000000111101011000101",
		b"00000000000111110111101010",
		b"00000000001000000011111001",
		b"00000000001000001111110011",
		b"00000000001000011011011000",
		b"00000000001000100110100110",
		b"00000000001000110001011111",
		b"00000000001000111100000010",
		b"00000000001001000110001101",
		b"00000000001001010000000010",
		b"00000000001001011001011111",
		b"00000000001001100010100110",
		b"00000000001001101011010100",
		b"00000000001001110011101011",
		b"00000000001001111011101001",
		b"00000000001010000011001111",
		b"00000000001010001010011101",
		b"00000000001010010001010011",
		b"00000000001010010111101111",
		b"00000000001010011101110011",
		b"00000000001010100011011101",
		b"00000000001010101000101111",
		b"00000000001010101101100111",
		b"00000000001010110010000110",
		b"00000000001010110110001100",
		b"00000000001010111001111000",
		b"00000000001010111101001011",
		b"00000000001011000000000100",
		b"00000000001011000010100100",
		b"00000000001011000100101011",
		b"00000000001011000110011000",
		b"00000000001011000111101011",
		b"00000000001011001000100101",
		b"00000000001011001001000110",
		b"00000000001011001001001101",
		b"00000000001011001000111011",
		b"00000000001011001000010000",
		b"00000000001011000111001100",
		b"00000000001011000101101111",
		b"00000000001011000011111001",
		b"00000000001011000001101011",
		b"00000000001010111111000100",
		b"00000000001010111100000101",
		b"00000000001010111000101101",
		b"00000000001010110100111110",
		b"00000000001010110000110110",
		b"00000000001010101100010111",
		b"00000000001010100111100001",
		b"00000000001010100010010100",
		b"00000000001010011100101111",
		b"00000000001010010110110100",
		b"00000000001010010000100011",
		b"00000000001010001001111011",
		b"00000000001010000010111110",
		b"00000000001001111011101011",
		b"00000000001001110100000011",
		b"00000000001001101100000110",
		b"00000000001001100011110101",
		b"00000000001001011011001111",
		b"00000000001001010010010101",
		b"00000000001001001001001000",
		b"00000000001000111111101000",
		b"00000000001000110101110100",
		b"00000000001000101011101110",
		b"00000000001000100001010111",
		b"00000000001000010110101101",
		b"00000000001000001011110010",
		b"00000000001000000000100111",
		b"00000000000111110101001010",
		b"00000000000111101001011110",
		b"00000000000111011101100010",
		b"00000000000111010001010111",
		b"00000000000111000100111110",
		b"00000000000110111000010110",
		b"00000000000110101011100000",
		b"00000000000110011110011101",
		b"00000000000110010001001100",
		b"00000000000110000011110000",
		b"00000000000101110110000111",
		b"00000000000101101000010011",
		b"00000000000101011010010100",
		b"00000000000101001100001010",
		b"00000000000100111101110110",
		b"00000000000100101111011001",
		b"00000000000100100000110011",
		b"00000000000100010010000100",
		b"00000000000100000011001101",
		b"00000000000011110100001110",
		b"00000000000011100101001001",
		b"00000000000011010101111100",
		b"00000000000011000110101010",
		b"00000000000010110111010010",
		b"00000000000010100111110101",
		b"00000000000010011000010100",
		b"00000000000010001000101111",
		b"00000000000001111001000110",
		b"00000000000001101001011010",
		b"00000000000001011001101011",
		b"00000000000001001001111011",
		b"00000000000000111010001001",
		b"00000000000000101010010110",
		b"00000000000000011010100011",
		b"00000000000000001010110000",
		b"11111111111111111010111101",
		b"11111111111111101011001100",
		b"11111111111111011011011100",
		b"11111111111111001011101110",
		b"11111111111110111100000010",
		b"11111111111110101100011010",
		b"11111111111110011100110101",
		b"11111111111110001101010100",
		b"11111111111101111101111000",
		b"11111111111101101110100000",
		b"11111111111101011111001110",
		b"11111111111101010000000010",
		b"11111111111101000000111101",
		b"11111111111100110001111110",
		b"11111111111100100011000110",
		b"11111111111100010100010110",
		b"11111111111100000101101110",
		b"11111111111011110111001111",
		b"11111111111011101000111001",
		b"11111111111011011010101100",
		b"11111111111011001100101001",
		b"11111111111010111110110001",
		b"11111111111010110001000011",
		b"11111111111010100011100000",
		b"11111111111010010110001001",
		b"11111111111010001000111101",
		b"11111111111001111011111110",
		b"11111111111001101111001011",
		b"11111111111001100010100110",
		b"11111111111001010110001101",
		b"11111111111001001010000011",
		b"11111111111000111110000110",
		b"11111111111000110010011000",
		b"11111111111000100110111000",
		b"11111111111000011011100111",
		b"11111111111000010000100110",
		b"11111111111000000101110100",
		b"11111111110111111011010001",
		b"11111111110111110001000000",
		b"11111111110111100110111110",
		b"11111111110111011101001101",
		b"11111111110111010011101101",
		b"11111111110111001010011110",
		b"11111111110111000001100000",
		b"11111111110110111000110101",
		b"11111111110110110000011010",
		b"11111111110110101000010010",
		b"11111111110110100000011100",
		b"11111111110110011000111001",
		b"11111111110110010001101000",
		b"11111111110110001010101010",
		b"11111111110110000011111110",
		b"11111111110101111101100110",
		b"11111111110101110111100001",
		b"11111111110101110001101111",
		b"11111111110101101100010000",
		b"11111111110101100111000101",
		b"11111111110101100010001110",
		b"11111111110101011101101010",
		b"11111111110101011001011010",
		b"11111111110101010101011101",
		b"11111111110101010001110101",
		b"11111111110101001110100001",
		b"11111111110101001011100000",
		b"11111111110101001000110011",
		b"11111111110101000110011011",
		b"11111111110101000100010110",
		b"11111111110101000010100101",
		b"11111111110101000001001001",
		b"11111111110101000000000000",
		b"11111111110100111111001011",
		b"11111111110100111110101010",
		b"11111111110100111110011100",
		b"11111111110100111110100011",
		b"11111111110100111110111101",
		b"11111111110100111111101010",
		b"11111111110101000000101011",
		b"11111111110101000010000000",
		b"11111111110101000011100111",
		b"11111111110101000101100010",
		b"11111111110101000111110000",
		b"11111111110101001010010001",
		b"11111111110101001101000100",
		b"11111111110101010000001010",
		b"11111111110101010011100010",
		b"11111111110101010111001100",
		b"11111111110101011011001001",
		b"11111111110101011111010111",
		b"11111111110101100011110111",
		b"11111111110101101000101001",
		b"11111111110101101101101011",
		b"11111111110101110010111111",
		b"11111111110101111000100011",
		b"11111111110101111110011000",
		b"11111111110110000100011101",
		b"11111111110110001010110010",
		b"11111111110110010001010111",
		b"11111111110110011000001100",
		b"11111111110110011111001111",
		b"11111111110110100110100010",
		b"11111111110110101110000011",
		b"11111111110110110101110011",
		b"11111111110110111101110000",
		b"11111111110111000101111100",
		b"11111111110111001110010101",
		b"11111111110111010110111011",
		b"11111111110111011111101101",
		b"11111111110111101000101101",
		b"11111111110111110001111000",
		b"11111111110111111011001111",
		b"11111111111000000100110010",
		b"11111111111000001110100000",
		b"11111111111000011000011001",
		b"11111111111000100010011100",
		b"11111111111000101100101001",
		b"11111111111000110110111111",
		b"11111111111001000001011111",
		b"11111111111001001100001001",
		b"11111111111001010110111010",
		b"11111111111001100001110100",
		b"11111111111001101100110110",
		b"11111111111001110111111111",
		b"11111111111010000011001111",
		b"11111111111010001110100110",
		b"11111111111010011010000011",
		b"11111111111010100101100110",
		b"11111111111010110001001111",
		b"11111111111010111100111100",
		b"11111111111011001000101111",
		b"11111111111011010100100110",
		b"11111111111011100000100000",
		b"11111111111011101100011110",
		b"11111111111011111000100000",
		b"11111111111100000100100100",
		b"11111111111100010000101010",
		b"11111111111100011100110010",
		b"11111111111100101000111100",
		b"11111111111100110101000111",
		b"11111111111101000001010011",
		b"11111111111101001101011111",
		b"11111111111101011001101011",
		b"11111111111101100101110111",
		b"11111111111101110010000001",
		b"11111111111101111110001011",
		b"11111111111110001010010011",
		b"11111111111110010110011001",
		b"11111111111110100010011100",
		b"11111111111110101110011101",
		b"11111111111110111010011010",
		b"11111111111111000110010100",
		b"11111111111111010010001010",
		b"11111111111111011101111100",
		b"11111111111111101001101001",
		b"11111111111111110101010001",
		b"00000000000000000000110100",
		b"00000000000000001100010001",
		b"00000000000000010111100111",
		b"00000000000000100010111000",
		b"00000000000000101110000001",
		b"00000000000000111001000100",
		b"00000000000001000011111110",
		b"00000000000001001110110001",
		b"00000000000001011001011100",
		b"00000000000001100011111110",
		b"00000000000001101110011000",
		b"00000000000001111000101000",
		b"00000000000010000010101111",
		b"00000000000010001100101100",
		b"00000000000010010110011111",
		b"00000000000010100000001000",
		b"00000000000010101001100110",
		b"00000000000010110010111001",
		b"00000000000010111100000001",
		b"00000000000011000100111101",
		b"00000000000011001101101110",
		b"00000000000011010110010011",
		b"00000000000011011110101011",
		b"00000000000011100110110111",
		b"00000000000011101110110110",
		b"00000000000011110110101000",
		b"00000000000011111110001101",
		b"00000000000100000101100100",
		b"00000000000100001100101110",
		b"00000000000100010011101010",
		b"00000000000100011010010111",
		b"00000000000100100000110111",
		b"00000000000100100111001000",
		b"00000000000100101101001010",
		b"00000000000100110010111101",
		b"00000000000100111000100010",
		b"00000000000100111101110111",
		b"00000000000101000010111101",
		b"00000000000101000111110100",
		b"00000000000101001100011011",
		b"00000000000101010000110010",
		b"00000000000101010100111001",
		b"00000000000101011000110001",
		b"00000000000101011100011000",
		b"00000000000101011111101111",
		b"00000000000101100010110110",
		b"00000000000101100101101101",
		b"00000000000101101000010011",
		b"00000000000101101010101001",
		b"00000000000101101100101110",
		b"00000000000101101110100010",
		b"00000000000101110000000110",
		b"00000000000101110001011001",
		b"00000000000101110010011011",
		b"00000000000101110011001100",
		b"00000000000101110011101101",
		b"00000000000101110011111101",
		b"00000000000101110011111100",
		b"00000000000101110011101010",
		b"00000000000101110011000111",
		b"00000000000101110010010100",
		b"00000000000101110001001111",
		b"00000000000101101111111010",
		b"00000000000101101110010101",
		b"00000000000101101100011110",
		b"00000000000101101010011000",
		b"00000000000101101000000000",
		b"00000000000101100101011000",
		b"00000000000101100010100000",
		b"00000000000101011111010111",
		b"00000000000101011011111110",
		b"00000000000101011000010101",
		b"00000000000101010100011100",
		b"00000000000101010000010011",
		b"00000000000101001011111010",
		b"00000000000101000111010010",
		b"00000000000101000010011010",
		b"00000000000100111101010010",
		b"00000000000100110111111100",
		b"00000000000100110010010110",
		b"00000000000100101100100001",
		b"00000000000100100110011101",
		b"00000000000100100000001011",
		b"00000000000100011001101010",
		b"00000000000100010010111010",
		b"00000000000100001011111101",
		b"00000000000100000100110010",
		b"00000000000011111101011000",
		b"00000000000011110101110010",
		b"00000000000011101101111110",
		b"00000000000011100101111100",
		b"00000000000011011101101110",
		b"00000000000011010101010011",
		b"00000000000011001100101011",
		b"00000000000011000011111000",
		b"00000000000010111010111000",
		b"00000000000010110001101100",
		b"00000000000010101000010101",
		b"00000000000010011110110010",
		b"00000000000010010101000100",
		b"00000000000010001011001100",
		b"00000000000010000001001000",
		b"00000000000001110110111011",
		b"00000000000001101100100011",
		b"00000000000001100010000010",
		b"00000000000001010111010111",
		b"00000000000001001100100011",
		b"00000000000001000001100101",
		b"00000000000000110110011111",
		b"00000000000000101011010001",
		b"00000000000000011111111010",
		b"00000000000000010100011100",
		b"00000000000000001000110110",
		b"11111111111111111101001000",
		b"11111111111111110001010100",
		b"11111111111111100101011001",
		b"11111111111111011001010111",
		b"11111111111111001101001111",
		b"11111111111111000001000010",
		b"11111111111110110100101111",
		b"11111111111110101000010110",
		b"11111111111110011011111001",
		b"11111111111110001111010111",
		b"11111111111110000010110001",
		b"11111111111101110110000111",
		b"11111111111101101001011001",
		b"11111111111101011100101000",
		b"11111111111101001111110100",
		b"11111111111101000010111100",
		b"11111111111100110110000011",
		b"11111111111100101001000111",
		b"11111111111100011100001001",
		b"11111111111100001111001010",
		b"11111111111100000010001001",
		b"11111111111011110101001000",
		b"11111111111011101000000110",
		b"11111111111011011011000011",
		b"11111111111011001110000000",
		b"11111111111011000000111110",
		b"11111111111010110011111100",
		b"11111111111010100110111011",
		b"11111111111010011001111100",
		b"11111111111010001100111101",
		b"11111111111010000000000001",
		b"11111111111001110011000110",
		b"11111111111001100110001110",
		b"11111111111001011001011001",
		b"11111111111001001100100110",
		b"11111111111000111111110110",
		b"11111111111000110011001010",
		b"11111111111000100110100010",
		b"11111111111000011001111110",
		b"11111111111000001101011110",
		b"11111111111000000001000011",
		b"11111111110111110100101100",
		b"11111111110111101000011011",
		b"11111111110111011100001111",
		b"11111111110111010000001000",
		b"11111111110111000100001000",
		b"11111111110110111000001110",
		b"11111111110110101100011010",
		b"11111111110110100000101101",
		b"11111111110110010101000110",
		b"11111111110110001001100111",
		b"11111111110101111110001111",
		b"11111111110101110010111111",
		b"11111111110101100111110111",
		b"11111111110101011100110111",
		b"11111111110101010001111111",
		b"11111111110101000111001111",
		b"11111111110100111100101001",
		b"11111111110100110010001011",
		b"11111111110100100111110110",
		b"11111111110100011101101011",
		b"11111111110100010011101001",
		b"11111111110100001001110001",
		b"11111111110100000000000011",
		b"11111111110011110110100000",
		b"11111111110011101101000110",
		b"11111111110011100011110111",
		b"11111111110011011010110010",
		b"11111111110011010001111001",
		b"11111111110011001001001010",
		b"11111111110011000000100110",
		b"11111111110010111000001110",
		b"11111111110010110000000001",
		b"11111111110010101000000000",
		b"11111111110010100000001010",
		b"11111111110010011000100000",
		b"11111111110010010001000011",
		b"11111111110010001001110001",
		b"11111111110010000010101100",
		b"11111111110001111011110010",
		b"11111111110001110101000110",
		b"11111111110001101110100110",
		b"11111111110001101000010010",
		b"11111111110001100010001011",
		b"11111111110001011100010001",
		b"11111111110001010110100100",
		b"11111111110001010001000100",
		b"11111111110001001011110001",
		b"11111111110001000110101011",
		b"11111111110001000001110011",
		b"11111111110000111101000111",
		b"11111111110000111000101001",
		b"11111111110000110100011000",
		b"11111111110000110000010101",
		b"11111111110000101100011111",
		b"11111111110000101000110110",
		b"11111111110000100101011011",
		b"11111111110000100010001110",
		b"11111111110000011111001110",
		b"11111111110000011100011100",
		b"11111111110000011001110111",
		b"11111111110000010111100000",
		b"11111111110000010101010110",
		b"11111111110000010011011010",
		b"11111111110000010001101100",
		b"11111111110000010000001011",
		b"11111111110000001110110111",
		b"11111111110000001101110001",
		b"11111111110000001100111001",
		b"11111111110000001100001110",
		b"11111111110000001011110001",
		b"11111111110000001011100000",
		b"11111111110000001011011101",
		b"11111111110000001011101000",
		b"11111111110000001100000000",
		b"11111111110000001100100100",
		b"11111111110000001101010110",
		b"11111111110000001110010101",
		b"11111111110000001111100001",
		b"11111111110000010000111010",
		b"11111111110000010010100000",
		b"11111111110000010100010010",
		b"11111111110000010110010001",
		b"11111111110000011000011100",
		b"11111111110000011010110100",
		b"11111111110000011101011001",
		b"11111111110000100000001001",
		b"11111111110000100011000110",
		b"11111111110000100110001111",
		b"11111111110000101001100100",
		b"11111111110000101101000100",
		b"11111111110000110000110001",
		b"11111111110000110100101001",
		b"11111111110000111000101100",
		b"11111111110000111100111011",
		b"11111111110001000001010100",
		b"11111111110001000101111001",
		b"11111111110001001010101001",
		b"11111111110001001111100100",
		b"11111111110001010100101001",
		b"11111111110001011001111001",
		b"11111111110001011111010011",
		b"11111111110001100100111000",
		b"11111111110001101010100110",
		b"11111111110001110000011110",
		b"11111111110001110110100000",
		b"11111111110001111100101100",
		b"11111111110010000011000001",
		b"11111111110010001001100000",
		b"11111111110010010000000111",
		b"11111111110010010110111000",
		b"11111111110010011101110001",
		b"11111111110010100100110011",
		b"11111111110010101011111101",
		b"11111111110010110011001111",
		b"11111111110010111010101010",
		b"11111111110011000010001100",
		b"11111111110011001001110110",
		b"11111111110011010001101000",
		b"11111111110011011001100001",
		b"11111111110011100001100001",
		b"11111111110011101001101000",
		b"11111111110011110001110110",
		b"11111111110011111010001011",
		b"11111111110100000010100110",
		b"11111111110100001011000111",
		b"11111111110100010011101111",
		b"11111111110100011100011100",
		b"11111111110100100101001111",
		b"11111111110100101110001000",
		b"11111111110100110111000101",
		b"11111111110101000000001000",
		b"11111111110101001001010000",
		b"11111111110101010010011101",
		b"11111111110101011011101110",
		b"11111111110101100101000100",
		b"11111111110101101110011101",
		b"11111111110101110111111011",
		b"11111111110110000001011101",
		b"11111111110110001011000010",
		b"11111111110110010100101010",
		b"11111111110110011110010110",
		b"11111111110110101000000101",
		b"11111111110110110001110111",
		b"11111111110110111011101011",
		b"11111111110111000101100010",
		b"11111111110111001111011011",
		b"11111111110111011001010111",
		b"11111111110111100011010100",
		b"11111111110111101101010011",
		b"11111111110111110111010100",
		b"11111111111000000001010110",
		b"11111111111000001011011001",
		b"11111111111000010101011101",
		b"11111111111000011111100010",
		b"11111111111000101001101000",
		b"11111111111000110011101110",
		b"11111111111000111101110101",
		b"11111111111001000111111100",
		b"11111111111001010010000010",
		b"11111111111001011100001001",
		b"11111111111001100110001111",
		b"11111111111001110000010101",
		b"11111111111001111010011010",
		b"11111111111010000100011110",
		b"11111111111010001110100001",
		b"11111111111010011000100011",
		b"11111111111010100010100100",
		b"11111111111010101100100011",
		b"11111111111010110110100001",
		b"11111111111011000000011101",
		b"11111111111011001010010111",
		b"11111111111011010100001110",
		b"11111111111011011110000100",
		b"11111111111011100111110111",
		b"11111111111011110001101000",
		b"11111111111011111011010110",
		b"11111111111100000101000001",
		b"11111111111100001110101010",
		b"11111111111100011000001111",
		b"11111111111100100001110001",
		b"11111111111100101011010000",
		b"11111111111100110100101011",
		b"11111111111100111110000011",
		b"11111111111101000111010111",
		b"11111111111101010000100111",
		b"11111111111101011001110011",
		b"11111111111101100010111100",
		b"11111111111101101100000000",
		b"11111111111101110101000000",
		b"11111111111101111101111011",
		b"11111111111110000110110010",
		b"11111111111110001111100101",
		b"11111111111110011000010010",
		b"11111111111110100000111011",
		b"11111111111110101001011111",
		b"11111111111110110001111111",
		b"11111111111110111010011001",
		b"11111111111111000010101110",
		b"11111111111111001010111101",
		b"11111111111111010011001000",
		b"11111111111111011011001101",
		b"11111111111111100011001100",
		b"11111111111111101011000110",
		b"11111111111111110010111010",
		b"11111111111111111010101001",
		b"00000000000000000010010010",
		b"00000000000000001001110101",
		b"00000000000000010001010010",
		b"00000000000000011000101010",
		b"00000000000000011111111011",
		b"00000000000000100111000110",
		b"00000000000000101110001011",
		b"00000000000000110101001010",
		b"00000000000000111100000011",
		b"00000000000001000010110101",
		b"00000000000001001001100001",
		b"00000000000001010000000111",
		b"00000000000001010110100111",
		b"00000000000001011101000000",
		b"00000000000001100011010010",
		b"00000000000001101001011110",
		b"00000000000001101111100100",
		b"00000000000001110101100011",
		b"00000000000001111011011100",
		b"00000000000010000001001110",
		b"00000000000010000110111001",
		b"00000000000010001100011110",
		b"00000000000010010001111100",
		b"00000000000010010111010100",
		b"00000000000010011100100101",
		b"00000000000010100001101111",
		b"00000000000010100110110011",
		b"00000000000010101011101111",
		b"00000000000010110000100110",
		b"00000000000010110101010101",
		b"00000000000010111001111110",
		b"00000000000010111110100001",
		b"00000000000011000010111100",
		b"00000000000011000111010001",
		b"00000000000011001011100000",
		b"00000000000011001111101000",
		b"00000000000011010011101001",
		b"00000000000011010111100100",
		b"00000000000011011011011000",
		b"00000000000011011111000101",
		b"00000000000011100010101100",
		b"00000000000011100110001101",
		b"00000000000011101001100111",
		b"00000000000011101100111010",
		b"00000000000011110000001000",
		b"00000000000011110011001111",
		b"00000000000011110110001111",
		b"00000000000011111001001001",
		b"00000000000011111011111101",
		b"00000000000011111110101011",
		b"00000000000100000001010010",
		b"00000000000100000011110011",
		b"00000000000100000110001111",
		b"00000000000100001000100100",
		b"00000000000100001010110011",
		b"00000000000100001100111100",
		b"00000000000100001110111111",
		b"00000000000100010000111100",
		b"00000000000100010010110100",
		b"00000000000100010100100101",
		b"00000000000100010110010001",
		b"00000000000100010111110111",
		b"00000000000100011001011000",
		b"00000000000100011010110011",
		b"00000000000100011100001000",
		b"00000000000100011101011000",
		b"00000000000100011110100010",
		b"00000000000100011111101000",
		b"00000000000100100000100111",
		b"00000000000100100001100010",
		b"00000000000100100010011000",
		b"00000000000100100011001000",
		b"00000000000100100011110011",
		b"00000000000100100100011010",
		b"00000000000100100100111011",
		b"00000000000100100101010111",
		b"00000000000100100101101111",
		b"00000000000100100110000010",
		b"00000000000100100110010001",
		b"00000000000100100110011010",
		b"00000000000100100110100000",
		b"00000000000100100110100001",
		b"00000000000100100110011101",
		b"00000000000100100110010101",
		b"00000000000100100110001001",
		b"00000000000100100101111001",
		b"00000000000100100101100100",
		b"00000000000100100101001100",
		b"00000000000100100100101111",
		b"00000000000100100100001111",
		b"00000000000100100011101011",
		b"00000000000100100011000011",
		b"00000000000100100010011000",
		b"00000000000100100001101000",
		b"00000000000100100000110110",
		b"00000000000100011111111111",
		b"00000000000100011111000110",
		b"00000000000100011110001001",
		b"00000000000100011101001001",
		b"00000000000100011100000101",
		b"00000000000100011010111111",
		b"00000000000100011001110101",
		b"00000000000100011000101001",
		b"00000000000100010111011010",
		b"00000000000100010110000111",
		b"00000000000100010100110011",
		b"00000000000100010011011011",
		b"00000000000100010010000001",
		b"00000000000100010000100100",
		b"00000000000100001111000101",
		b"00000000000100001101100011",
		b"00000000000100001011111111",
		b"00000000000100001010011001",
		b"00000000000100001000110000",
		b"00000000000100000111000110",
		b"00000000000100000101011001",
		b"00000000000100000011101010",
		b"00000000000100000001111010",
		b"00000000000100000000000111",
		b"00000000000011111110010011",
		b"00000000000011111100011101",
		b"00000000000011111010100101",
		b"00000000000011111000101100",
		b"00000000000011110110110001",
		b"00000000000011110100110101",
		b"00000000000011110010110111",
		b"00000000000011110000111000",
		b"00000000000011101110110111",
		b"00000000000011101100110110",
		b"00000000000011101010110011",
		b"00000000000011101000101111",
		b"00000000000011100110101010",
		b"00000000000011100100100100",
		b"00000000000011100010011101",
		b"00000000000011100000010110",
		b"00000000000011011110001101",
		b"00000000000011011100000100",
		b"00000000000011011001111001",
		b"00000000000011010111101111",
		b"00000000000011010101100011",
		b"00000000000011010011010111",
		b"00000000000011010001001011",
		b"00000000000011001110111110",
		b"00000000000011001100110001",
		b"00000000000011001010100011",
		b"00000000000011001000010101",
		b"00000000000011000110000111",
		b"00000000000011000011111000",
		b"00000000000011000001101010",
		b"00000000000010111111011011",
		b"00000000000010111101001100",
		b"00000000000010111010111101",
		b"00000000000010111000101111",
		b"00000000000010110110100000",
		b"00000000000010110100010001",
		b"00000000000010110010000011",
		b"00000000000010101111110100",
		b"00000000000010101101100110",
		b"00000000000010101011011000",
		b"00000000000010101001001011",
		b"00000000000010100110111101",
		b"00000000000010100100110000",
		b"00000000000010100010100100",
		b"00000000000010100000011000",
		b"00000000000010011110001100",
		b"00000000000010011100000001",
		b"00000000000010011001110110",
		b"00000000000010010111101100",
		b"00000000000010010101100011",
		b"00000000000010010011011010",
		b"00000000000010010001010010",
		b"00000000000010001111001010",
		b"00000000000010001101000100",
		b"00000000000010001010111110",
		b"00000000000010001000111000",
		b"00000000000010000110110100",
		b"00000000000010000100110000",
		b"00000000000010000010101101",
		b"00000000000010000000101011",
		b"00000000000001111110101010",
		b"00000000000001111100101010",
		b"00000000000001111010101010",
		b"00000000000001111000101100",
		b"00000000000001110110101110",
		b"00000000000001110100110010",
		b"00000000000001110010110110",
		b"00000000000001110000111100",
		b"00000000000001101111000010",
		b"00000000000001101101001010",
		b"00000000000001101011010011",
		b"00000000000001101001011100",
		b"00000000000001100111100111",
		b"00000000000001100101110011",
		b"00000000000001100100000000",
		b"00000000000001100010001110",
		b"00000000000001100000011101",
		b"00000000000001011110101101",
		b"00000000000001011100111111",
		b"00000000000001011011010001",
		b"00000000000001011001100101",
		b"00000000000001010111111010",
		b"00000000000001010110010000",
		b"00000000000001010100100111",
		b"00000000000001010011000000",
		b"00000000000001010001011010",
		b"00000000000001001111110100",
		b"00000000000001001110010000",
		b"00000000000001001100101110",
		b"00000000000001001011001100",
		b"00000000000001001001101100",
		b"00000000000001001000001101",
		b"00000000000001000110101111",
		b"00000000000001000101010010",
		b"00000000000001000011110111",
		b"00000000000001000010011101",
		b"00000000000001000001000100",
		b"00000000000000111111101100",
		b"00000000000000111110010101",
		b"00000000000000111101000000",
		b"00000000000000111011101100",
		b"00000000000000111010011001",
		b"00000000000000111001000111",
		b"00000000000000110111110111",
		b"00000000000000110110100111",
		b"00000000000000110101011001",
		b"00000000000000110100001100",
		b"00000000000000110011000000",
		b"00000000000000110001110110",
		b"00000000000000110000101100",
		b"00000000000000101111100100",
		b"00000000000000101110011101",
		b"00000000000000101101010111",
		b"00000000000000101100010010",
		b"00000000000000101011001111",
		b"00000000000000101010001100",
		b"00000000000000101001001011",
		b"00000000000000101000001011",
		b"00000000000000100111001100",
		b"00000000000000100110001110",
		b"00000000000000100101010001",
		b"00000000000000100100010101",
		b"00000000000000100011011010",
		b"00000000000000100010100001",
		b"00000000000000100001101000",
		b"00000000000000100000110001",
		b"00000000000000011111111010",
		b"00000000000000011111000101",
		b"00000000000000011110010000",
		b"00000000000000011101011101",
		b"00000000000000011100101010",
		b"00000000000000011011111001",
		b"00000000000000011011001001",
		b"00000000000000011010011001",
		b"00000000000000011001101011",
		b"00000000000000011000111101",
		b"00000000000000011000010001",
		b"00000000000000010111100101",
		b"00000000000000010110111010",
		b"00000000000000010110010000",
		b"00000000000000010101100111",
		b"00000000000000010100111111",
		b"00000000000000010100011000",
		b"00000000000000010011110010",
		b"00000000000000010011001100",
		b"00000000000000010010101000",
		b"00000000000000010010000100",
		b"00000000000000010001100001",
		b"00000000000000010000111111",
		b"00000000000000010000011110",
		b"00000000000000001111111101",
		b"00000000000000001111011101",
		b"00000000000000001110111110",
		b"00000000000000001110100000",
		b"00000000000000001110000010",
		b"00000000000000001101100101",
		b"00000000000000001101001001",
		b"00000000000000001100101110",
		b"00000000000000001100010011",
		b"00000000000000001011111001",
		b"00000000000000001011100000",
		b"00000000000000001011000111",
		b"00000000000000001010101111",
		b"00000000000000001010010111",
		b"00000000000000001010000001",
		b"00000000000000001001101010",
		b"00000000000000001001010101",
		b"00000000000000001001000000",
		b"00000000000000001000101011",
		b"00000000000000001000010111",
		b"00000000000000001000000100",
		b"00000000000000000111110001",
		b"00000000000000000111011111",
		b"00000000000000000111001101",
		b"00000000000000000110111100",
		b"00000000000000000110101011",
		b"00000000000000000110011011",
		b"00000000000000000110001011",
		b"00000000000000000101111100",
		b"00000000000000000101101101",
		b"00000000000000000101011111",
		b"00000000000000000101010001",
		b"00000000000000000101000100",
		b"00000000000000000100110110",
		b"00000000000000000100101010",
		b"00000000000000000100011110",
		b"00000000000000000100010010",
		b"00000000000000000100000110",
		b"00000000000000000011111011",
		b"00000000000000000011110000",
		b"00000000000000000011100110",
		b"00000000000000000011011100",
		b"00000000000000000011010010",
		b"00000000000000000011001001",
		b"00000000000000000011000000",
		b"00000000000000000010110111",
		b"00000000000000000010101111",
		b"00000000000000000010100111",
		b"00000000000000000010011111",
		b"00000000000000000010011000",
		b"00000000000000000010010000",
		b"00000000000000000010001010",
		b"00000000000000000010000011",
		b"00000000000000000001111100",
		b"00000000000000000001110110",
		b"00000000000000000001110000",
		b"00000000000000000001101011",
		b"00000000000000000001100101",
		b"00000000000000000001100000",
		b"00000000000000000001011011",
		b"00000000000000000001010110",
		b"00000000000000000001010001",
		b"00000000000000000001001101",
		b"00000000000000000001001000",
		b"00000000000000000001000100",
		b"00000000000000000001000000",
		b"00000000000000000000111101",
		b"00000000000000000000111001",
		b"00000000000000000000110110",
		b"00000000000000000000110010",
		b"00000000000000000000101111",
		b"00000000000000000000101100",
		b"00000000000000000000101010",
		b"00000000000000000000100111",
		b"00000000000000000000100100",
		b"00000000000000000000100010",
		b"00000000000000000000100000",
		b"00000000000000000000011101",
		b"00000000000000000000011011",
		b"00000000000000000000011001",
		b"00000000000000000000010111",
		b"00000000000000000000010110",
		b"00000000000000000000010100",
		b"00000000000000000000010010",
		b"00000000000000000000010001",
		b"00000000000000000000001111",
		b"00000000000000000000001110",
		b"00000000000000000000001101",
		b"00000000000000000000001100",
		b"00000000000000000000001011",
		b"00000000000000000000001010",
		b"00000000000000000000001001",
		b"00000000000000000000001000",
		b"00000000000000000000000111",
		b"00000000000000000000000110",
		b"00000000000000000000000101",
		b"00000000000000000000000101",
		b"00000000000000000000000100",
		b"00000000000000000000000100",
		b"00000000000000000000000011",
		b"00000000000000000000000011",
		b"00000000000000000000000010",
		b"00000000000000000000000010",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"11111111111111111111111111",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000001",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000",
		b"00000000000000000000000000"
	);

end src_rom_pkg;