library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package src_rom_pkg is

	constant COE_WIDTH	: integer := 24;
	constant COE_CENTRE	: signed( 23 downto 0 ) := b"011111110101110000101001";

	type COE_ROM_TYPE is array( 4095 downto 0 ) of signed( 23 downto 0 );
	constant COE_ROM	 : COE_ROM_TYPE := (
		b"011111110101100100011100",
		b"011111110100111111110100",
		b"011111110100000010110011",
		b"011111110010101101011010",
		b"011111110000111111101011",
		b"011111101110111001100111",
		b"011111101100011011010011",
		b"011111101001100100110001",
		b"011111100110010110000110",
		b"011111100010101111010101",
		b"011111011110110000100100",
		b"011111011010011001111001",
		b"011111010101101011011001",
		b"011111010000100101001010",
		b"011111001011000111010101",
		b"011111000101010010000000",
		b"011110111111000101010100",
		b"011110111000100001011000",
		b"011110110001100110010111",
		b"011110101010010100011010",
		b"011110100010101011101010",
		b"011110011010101100010011",
		b"011110010010010110011111",
		b"011110001001101010011001",
		b"011110000000101000001111",
		b"011101110111010000001011",
		b"011101101101100010011100",
		b"011101100011011111001110",
		b"011101011001000110101111",
		b"011101001110011001001101",
		b"011101000011010110111000",
		b"011100110111111111111110",
		b"011100101100010100101111",
		b"011100100000010101011010",
		b"011100010100000010010001",
		b"011100000111011011100100",
		b"011011111010100001100100",
		b"011011101101010100100010",
		b"011011011111110100110010",
		b"011011010010000010100101",
		b"011011000011111110001101",
		b"011010110101100111111111",
		b"011010100111000000001101",
		b"011010011000000111001011",
		b"011010001000111101001110",
		b"011001111001100010101010",
		b"011001101001110111110100",
		b"011001011001111101000001",
		b"011001001001110010100110",
		b"011000111001011000111010",
		b"011000101000110000010010",
		b"011000010111111001000100",
		b"011000000110110011101000",
		b"010111110101100000010100",
		b"010111100011111111100000",
		b"010111010010010001100010",
		b"010111000000010110110010",
		b"010110101110001111101001",
		b"010110011011111100011110",
		b"010110001001011101101010",
		b"010101110110110011100101",
		b"010101100011111110101000",
		b"010101010000111111001011",
		b"010100111101110101101001",
		b"010100101010100010011001",
		b"010100010111000101110110",
		b"010100000011100000011000",
		b"010011101111110010011010",
		b"010011011011111100010110",
		b"010011000111111110100100",
		b"010010110011111001100000",
		b"010010011111101101100011",
		b"010010001011011011001000",
		b"010001110111000010101000",
		b"010001100010100100011110",
		b"010001001110000001000100",
		b"010000111001011000110101",
		b"010000100100101100001011",
		b"010000001111111011100000",
		b"001111111011000111010000",
		b"001111100110001111110100",
		b"001111010001010101100111",
		b"001110111100011001000011",
		b"001110100111011010100011",
		b"001110010010011010100000",
		b"001101111101011001010111",
		b"001101101000010111100000",
		b"001101010011010101010110",
		b"001100111110010011010010",
		b"001100101001010001110000",
		b"001100010100010001001000",
		b"001011111111010001110101",
		b"001011101010010100010001",
		b"001011010101011000110100",
		b"001011000000011111111001",
		b"001010101011101001111000",
		b"001010010110110111001011",
		b"001010000010001000001011",
		b"001001101101011101001111",
		b"001001011000110110110010",
		b"001001000100010101001100",
		b"001000101111111000110100",
		b"001000011011100010000011",
		b"001000000111010001010000",
		b"000111110011000110110011",
		b"000111011111000011000011",
		b"000111001011000110010111",
		b"000110110111010001000111",
		b"000110100011100011101000",
		b"000110001111111110010001",
		b"000101111100100001011000",
		b"000101101001001101010010",
		b"000101010110000010010101",
		b"000101000011000000110111",
		b"000100110000001001001011",
		b"000100011101011011100111",
		b"000100001010111000011110",
		b"000011111000100000000101",
		b"000011100110010010101111",
		b"000011010100010000101111",
		b"000011000010011010010111",
		b"000010110000101111111011",
		b"000010011111010001101100",
		b"000010001101111111111101",
		b"000001111100111010111110",
		b"000001101100000011000000",
		b"000001011011011000010101",
		b"000001001010111011001011",
		b"000000111010101011110101",
		b"000000101010101010011111",
		b"000000011010110111011010",
		b"000000001011010010110011",
		b"111111111011111100111010",
		b"111111101100110101111100",
		b"111111011101111110000111",
		b"111111001111010101100110",
		b"111111000000111100101000",
		b"111110110010110011010111",
		b"111110100100111001111111",
		b"111110010111010000101101",
		b"111110001001110111101001",
		b"111101111100101110111111",
		b"111101101111110110111000",
		b"111101100011001111011111",
		b"111101010110111000111011",
		b"111101001010110011010101",
		b"111100111110111110110101",
		b"111100110011011011100100",
		b"111100101000001001100111",
		b"111100011101001001000110",
		b"111100010010011010000111",
		b"111100000111111100110000",
		b"111011111101110001000101",
		b"111011110011110111001100",
		b"111011101010001111001010",
		b"111011100000111001000001",
		b"111011010111110100110101",
		b"111011001111000010101010",
		b"111011000110100010100010",
		b"111010111110010100011110",
		b"111010110110011000100010",
		b"111010101110101110101101",
		b"111010100111010111000000",
		b"111010100000010001011100",
		b"111010011001011110000000",
		b"111010010010111100101100",
		b"111010001100101101011111",
		b"111010000110110000010110",
		b"111010000001000101010001",
		b"111001111011101100001100",
		b"111001110110100101000101",
		b"111001110001101111111000",
		b"111001101101001100100010",
		b"111001101000111010111110",
		b"111001100100111011001001",
		b"111001100001001100111100",
		b"111001011101110000010010",
		b"111001011010100101000110",
		b"111001010111101011010001",
		b"111001010101000010101101",
		b"111001010010101011010010",
		b"111001010000100100111001",
		b"111001001110101111011011",
		b"111001001101001010101111",
		b"111001001011110110101100",
		b"111001001010110011001010",
		b"111001001001111111111110",
		b"111001001001011101000001",
		b"111001001001001010000110",
		b"111001001001000111000101",
		b"111001001001010011110001",
		b"111001001001110000000000",
		b"111001001010011011101000",
		b"111001001011010110011011",
		b"111001001100100000001110",
		b"111001001101111000110101",
		b"111001001111100000000010",
		b"111001010001010101101000",
		b"111001010011011001011100",
		b"111001010101101011001110",
		b"111001011000001010110001",
		b"111001011010110111110111",
		b"111001011101110010010001",
		b"111001100000111001110010",
		b"111001100100001110001001",
		b"111001100111101111001000",
		b"111001101011011100100000",
		b"111001101111010110000000",
		b"111001110011011011011010",
		b"111001110111101100011101",
		b"111001111100001000111001",
		b"111010000000110000011101",
		b"111010000101100010111001",
		b"111010001010011111111100",
		b"111010001111100111010101",
		b"111010010100111000110011",
		b"111010011010010100000101",
		b"111010011111111000111001",
		b"111010100101100110111111",
		b"111010101011011110000011",
		b"111010110001011101110101",
		b"111010110111100110000010",
		b"111010111101110110011001",
		b"111011000100001110100111",
		b"111011001010101110011011",
		b"111011010001010101100010",
		b"111011011000000011101001",
		b"111011011110111000011111",
		b"111011100101110011110000",
		b"111011101100110101001011",
		b"111011110011111100011100",
		b"111011111011001001010010",
		b"111100000010011011011010",
		b"111100001001110010100000",
		b"111100010001001110010100",
		b"111100011000101110100001",
		b"111100100000010010110110",
		b"111100100111111011000000",
		b"111100101111100110101100",
		b"111100110111010101101000",
		b"111100111111000111100010",
		b"111101000110111100000111",
		b"111101001110110011000101",
		b"111101010110101100001010",
		b"111101011110100111000011",
		b"111101100110100011011110",
		b"111101101110100001001010",
		b"111101110110011111110101",
		b"111101111110011111001100",
		b"111110000110011110111111",
		b"111110001110011110111011",
		b"111110010110011110110000",
		b"111110011110011110001011",
		b"111110100110011100111101",
		b"111110101110011010110100",
		b"111110110110010111011110",
		b"111110111110010010101101",
		b"111111000110001100001110",
		b"111111001110000011110010",
		b"111111010101111001001001",
		b"111111011101101100000011",
		b"111111100101011100001111",
		b"111111101101001001100000",
		b"111111110100110011100100",
		b"111111111100011010001110",
		b"000000000011111101001110",
		b"000000001011011100010110",
		b"000000010010110111011000",
		b"000000011010001110000100",
		b"000000100001100000001110",
		b"000000101000101101100111",
		b"000000101111110110000010",
		b"000000110110111001010011",
		b"000000111101110111001011",
		b"000001000100101111011111",
		b"000001001011100010000010",
		b"000001010010001110101000",
		b"000001011000110101000101",
		b"000001011111010101001110",
		b"000001100101101110110111",
		b"000001101100000001110110",
		b"000001110010001110000000",
		b"000001111000010011001010",
		b"000001111110010001001010",
		b"000010000100000111111000",
		b"000010001001110111001000",
		b"000010001111011110110011",
		b"000010010100111110101110",
		b"000010011010010110110011",
		b"000010011111100110111000",
		b"000010100100101110110110",
		b"000010101001101110100100",
		b"000010101110100101111101",
		b"000010110011010100111001",
		b"000010110111111011010001",
		b"000010111100011000111111",
		b"000011000000101101111101",
		b"000011000100111010000110",
		b"000011001000111101010100",
		b"000011001100110111100010",
		b"000011010000101000101101",
		b"000011010100010000101110",
		b"000011010111101111100011",
		b"000011011011000101001000",
		b"000011011110010001011001",
		b"000011100001010100010100",
		b"000011100100001101110101",
		b"000011100110111101111011",
		b"000011101001100100100100",
		b"000011101100000001101110",
		b"000011101110010101010111",
		b"000011110000011111011111",
		b"000011110010100000000100",
		b"000011110100010111001000",
		b"000011110110000100101000",
		b"000011110111101000100110",
		b"000011111001000011000011",
		b"000011111010010011111110",
		b"000011111011011011011011",
		b"000011111100011001011001",
		b"000011111101001101111010",
		b"000011111101111001000010",
		b"000011111110011010110001",
		b"000011111110110011001100",
		b"000011111111000010010101",
		b"000011111111001000001111",
		b"000011111111000100111110",
		b"000011111110111000100110",
		b"000011111110100011001011",
		b"000011111110000100110001",
		b"000011111101011101011101",
		b"000011111100101101010101",
		b"000011111011110100011100",
		b"000011111010110010111010",
		b"000011111001101000110011",
		b"000011111000010110001110",
		b"000011110110111011010000",
		b"000011110101011000000001",
		b"000011110011101100100111",
		b"000011110001111001001010",
		b"000011101111111101101111",
		b"000011101101111010100000",
		b"000011101011101111100011",
		b"000011101001011101000000",
		b"000011100111000010111111",
		b"000011100100100001101001",
		b"000011100001111001000111",
		b"000011011111001001100000",
		b"000011011100010010111110",
		b"000011011001010101101001",
		b"000011010110010001101011",
		b"000011010011000111001110",
		b"000011001111110110011010",
		b"000011001100011111011011",
		b"000011001001000010011000",
		b"000011000101011111011101",
		b"000011000001110110110100",
		b"000010111110001000100110",
		b"000010111010010100111111",
		b"000010110110011100001001",
		b"000010110010011110001110",
		b"000010101110011011011001",
		b"000010101010010011110110",
		b"000010100110000111101110",
		b"000010100001110111001110",
		b"000010011101100010100000",
		b"000010011001001001110000",
		b"000010010100101101001000",
		b"000010010000001100110101",
		b"000010001011101001000010",
		b"000010000111000001111001",
		b"000010000010010111100111",
		b"000001111101101010011000",
		b"000001111000111010010110",
		b"000001110100000111101110",
		b"000001101111010010101011",
		b"000001101010011011011001",
		b"000001100101100010000011",
		b"000001100000100110110110",
		b"000001011011101001111101",
		b"000001010110101011100011",
		b"000001010001101011110101",
		b"000001001100101010111110",
		b"000001000111101001001001",
		b"000001000010100110100011",
		b"000000111101100011010111",
		b"000000111000011111110000",
		b"000000110011011011111001",
		b"000000101110010111111111",
		b"000000101001010100001101",
		b"000000100100010000101110",
		b"000000011111001101101101",
		b"000000011010001011010101",
		b"000000010101001001110010",
		b"000000010000001001001110",
		b"000000001011001001110100",
		b"000000000110001011101111",
		b"000000000001001111001011",
		b"111111111100010100010000",
		b"111111110111011011001011",
		b"111111110010100100000101",
		b"111111101101101111001000",
		b"111111101000111100011110",
		b"111111100100001100010011",
		b"111111011111011110101110",
		b"111111011010110011111011",
		b"111111010110001100000010",
		b"111111010001100111001101",
		b"111111001101000101100110",
		b"111111001000100111010101",
		b"111111000100001100100011",
		b"111110111111110101011001",
		b"111110111011100010000000",
		b"111110110111010010011111",
		b"111110110011000111000000",
		b"111110101110111111101011",
		b"111110101010111100100110",
		b"111110100110111101111011",
		b"111110100011000011110000",
		b"111110011111001110001100",
		b"111110011011011101011000",
		b"111110010111110001011001",
		b"111110010100001010010111",
		b"111110010000101000010111",
		b"111110001101001011100001",
		b"111110001001110011111010",
		b"111110000110100001101000",
		b"111110000011010100110001",
		b"111110000000001101011011",
		b"111101111101001011101001",
		b"111101111010001111100011",
		b"111101110111011001001100",
		b"111101110100101000101000",
		b"111101110001111101111101",
		b"111101101111011001001111",
		b"111101101100111010100000",
		b"111101101010100001110110",
		b"111101101000001111010010",
		b"111101100110000010111010",
		b"111101100011111100101111",
		b"111101100001111100110100",
		b"111101100000000011001101",
		b"111101011110001111111010",
		b"111101011100100010111110",
		b"111101011010111100011100",
		b"111101011001011100010100",
		b"111101011000000010101000",
		b"111101010110101111011010",
		b"111101010101100010101001",
		b"111101010100011100010111",
		b"111101010011011100100101",
		b"111101010010100011010010",
		b"111101010001110000011110",
		b"111101010001000100001010",
		b"111101010000011110010100",
		b"111101001111111110111100",
		b"111101001111100110000010",
		b"111101001111010011100100",
		b"111101001111000111100000",
		b"111101001111000001110110",
		b"111101001111000010100100",
		b"111101001111001001100110",
		b"111101001111010110111101",
		b"111101001111101010100100",
		b"111101010000000100011001",
		b"111101010000100100011010",
		b"111101010001001010100100",
		b"111101010001110110110011",
		b"111101010010101001000100",
		b"111101010011100001010011",
		b"111101010100011111011101",
		b"111101010101100011011101",
		b"111101010110101101010000",
		b"111101010111111100110001",
		b"111101011001010001111100",
		b"111101011010101100101100",
		b"111101011100001100111011",
		b"111101011101110010100110",
		b"111101011111011101100110",
		b"111101100001001101110111",
		b"111101100011000011010010",
		b"111101100100111101110011",
		b"111101100110111101010100",
		b"111101101001000001101101",
		b"111101101011001010111011",
		b"111101101101011000110101",
		b"111101101111101011010110",
		b"111101110010000010010110",
		b"111101110100011101110001",
		b"111101110110111101011110",
		b"111101111001100001010111",
		b"111101111100001001010101",
		b"111101111110110101010000",
		b"111110000001100101000010",
		b"111110000100011000100011",
		b"111110000111001111101100",
		b"111110001010001010010101",
		b"111110001101001000010110",
		b"111110010000001001101001",
		b"111110010011001110000100",
		b"111110010110010101100001",
		b"111110011001011111110111",
		b"111110011100101100111110",
		b"111110011111111100101111",
		b"111110100011001111000001",
		b"111110100110100011101100",
		b"111110101001111010101000",
		b"111110101101010011101100",
		b"111110110000101110110001",
		b"111110110100001011101110",
		b"111110110111101010011010",
		b"111110111011001010101101",
		b"111110111110101100100000",
		b"111111000010001111101001",
		b"111111000101110100000000",
		b"111111001001011001011100",
		b"111111001100111111110110",
		b"111111010000100111000100",
		b"111111010100001110111111",
		b"111111010111110111011110",
		b"111111011011100000011000",
		b"111111011111001001100110",
		b"111111100010110010111110",
		b"111111100110011100011001",
		b"111111101010000101101110",
		b"111111101101101110110101",
		b"111111110001010111100110",
		b"111111110100111111111000",
		b"111111111000100111100100",
		b"111111111100001110100010",
		b"111111111111110100101001",
		b"000000000011011001110010",
		b"000000000110111101110100",
		b"000000001010100000101001",
		b"000000001110000010000111",
		b"000000010001100010001001",
		b"000000010101000000100101",
		b"000000011000011101010101",
		b"000000011011111000010010",
		b"000000011111010001010011",
		b"000000100010101000010010",
		b"000000100101111101001000",
		b"000000101001001111101110",
		b"000000101100011111111100",
		b"000000101111101101101101",
		b"000000110010111000111010",
		b"000000110110000001011011",
		b"000000111001000111001011",
		b"000000111100001010000011",
		b"000000111111001001111110",
		b"000001000010000110110100",
		b"000001000101000000100001",
		b"000001000111110110111111",
		b"000001001010101010001000",
		b"000001001101011001110110",
		b"000001010000000110000100",
		b"000001010010101110101101",
		b"000001010101010011101100",
		b"000001010111110100111100",
		b"000001011010010010011000",
		b"000001011100101011111100",
		b"000001011111000001100100",
		b"000001100001010011001010",
		b"000001100011100000101011",
		b"000001100101101010000011",
		b"000001100111101111001111",
		b"000001101001110000001010",
		b"000001101011101100110000",
		b"000001101101100101000000",
		b"000001101111011000110101",
		b"000001110001001000001101",
		b"000001110010110011000101",
		b"000001110100011001011010",
		b"000001110101111011001001",
		b"000001110111011000010001",
		b"000001111000110000110000",
		b"000001111010000100100011",
		b"000001111011010011101000",
		b"000001111100011101111111",
		b"000001111101100011100101",
		b"000001111110100100011010",
		b"000001111111100000011011",
		b"000010000000010111101010",
		b"000010000001001010000011",
		b"000010000001110111101000",
		b"000010000010100000011000",
		b"000010000011000100010010",
		b"000010000011100011010110",
		b"000010000011111101100101",
		b"000010000100010010111111",
		b"000010000100100011100100",
		b"000010000100101111010110",
		b"000010000100110110010011",
		b"000010000100111000011111",
		b"000010000100110101111001",
		b"000010000100101110100100",
		b"000010000100100010100000",
		b"000010000100010001101111",
		b"000010000011111100010011",
		b"000010000011100010001110",
		b"000010000011000011100010",
		b"000010000010100000010001",
		b"000010000001111000011110",
		b"000010000001001100001011",
		b"000010000000011011011010",
		b"000001111111100110010000",
		b"000001111110101100101110",
		b"000001111101101110111000",
		b"000001111100101100110001",
		b"000001111011100110011100",
		b"000001111010011011111101",
		b"000001111001001101011001",
		b"000001110111111010110001",
		b"000001110110100100001011",
		b"000001110101001001101010",
		b"000001110011101011010100",
		b"000001110010001001001011",
		b"000001110000100011010100",
		b"000001101110111001110100",
		b"000001101101001100110000",
		b"000001101011011100001100",
		b"000001101001101000001101",
		b"000001100111110000111001",
		b"000001100101110110010011",
		b"000001100011111000100010",
		b"000001100001110111101010",
		b"000001011111110011110001",
		b"000001011101101100111101",
		b"000001011011100011010010",
		b"000001011001010110110111",
		b"000001010111000111110000",
		b"000001010100110110000101",
		b"000001010010100001111010",
		b"000001010000001011010101",
		b"000001001101110010011101",
		b"000001001011010111011000",
		b"000001001000111010001010",
		b"000001000110011010111100",
		b"000001000011111001110001",
		b"000001000001010110110010",
		b"000000111110110010000100",
		b"000000111100001011101101",
		b"000000111001100011110100",
		b"000000110110111010011111",
		b"000000110100001111110100",
		b"000000110001100011111011",
		b"000000101110110110111000",
		b"000000101100001000110011",
		b"000000101001011001110010",
		b"000000100110101001111011",
		b"000000100011111001010101",
		b"000000100001001000000111",
		b"000000011110010110010111",
		b"000000011011100100001011",
		b"000000011000110001101001",
		b"000000010101111110111001",
		b"000000010011001100000001",
		b"000000010000011001000110",
		b"000000001101100110010000",
		b"000000001010110011100100",
		b"000000001000000001001010",
		b"000000000101001111000111",
		b"000000000010011101100001",
		b"111111111111101100011111",
		b"111111111100111100001000",
		b"111111111010001100100000",
		b"111111110111011101101110",
		b"111111110100101111111001",
		b"111111110010000011000101",
		b"111111101111010111011010",
		b"111111101100101100111101",
		b"111111101010000011110011",
		b"111111100111011100000011",
		b"111111100100110101110001",
		b"111111100010010001000101",
		b"111111011111101110000010",
		b"111111011101001100101111",
		b"111111011010101101010001",
		b"111111011000001111101101",
		b"111111010101110100001000",
		b"111111010011011010101000",
		b"111111010001000011010001",
		b"111111001110101110001000",
		b"111111001100011011010011",
		b"111111001010001010110101",
		b"111111000111111100110011",
		b"111111000101110001010011",
		b"111111000011101000010111",
		b"111111000001100010000101",
		b"111110111111011110100001",
		b"111110111101011101101111",
		b"111110111011011111110010",
		b"111110111001100100101111",
		b"111110110111101100101010",
		b"111110110101110111100101",
		b"111110110100000101100100",
		b"111110110010010110101100",
		b"111110110000101010111110",
		b"111110101111000010011111",
		b"111110101101011101010000",
		b"111110101011111011010110",
		b"111110101010011100110010",
		b"111110101001000001100111",
		b"111110100111101001111001",
		b"111110100110010101101000",
		b"111110100101000100111000",
		b"111110100011110111101011",
		b"111110100010101110000001",
		b"111110100001100111111110",
		b"111110100000100101100011",
		b"111110011111100110110010",
		b"111110011110101011101011",
		b"111110011101110100010001",
		b"111110011101000000100011",
		b"111110011100010000100101",
		b"111110011011100100010101",
		b"111110011010111011110101",
		b"111110011010010111000110",
		b"111110011001110110001000",
		b"111110011001011000111100",
		b"111110011000111111100001",
		b"111110011000101001111000",
		b"111110011000011000000000",
		b"111110011000001001111010",
		b"111110010111111111100100",
		b"111110010111111001000000",
		b"111110010111110110001011",
		b"111110010111110111000110",
		b"111110010111111011101111",
		b"111110011000000100000101",
		b"111110011000010000001000",
		b"111110011000011111110110",
		b"111110011000110011001110",
		b"111110011001001010001101",
		b"111110011001100100110100",
		b"111110011010000010111111",
		b"111110011010100100101101",
		b"111110011011001001111101",
		b"111110011011110010101011",
		b"111110011100011110110110",
		b"111110011101001110011011",
		b"111110011110000001011001",
		b"111110011110110111101011",
		b"111110011111110001010001",
		b"111110100000101110000110",
		b"111110100001101110001001",
		b"111110100010110001010101",
		b"111110100011110111101001",
		b"111110100101000001000000",
		b"111110100110001101011000",
		b"111110100111011100101110",
		b"111110101000101110111101",
		b"111110101010000100000010",
		b"111110101011011011111001",
		b"111110101100110110100000",
		b"111110101110010011110001",
		b"111110101111110011101010",
		b"111110110001010110000110",
		b"111110110010111011000000",
		b"111110110100100010010110",
		b"111110110110001100000010",
		b"111110110111111000000001",
		b"111110111001100110001101",
		b"111110111011010110100100",
		b"111110111101001001000000",
		b"111110111110111101011100",
		b"111111000000110011110100",
		b"111111000010101100000100",
		b"111111000100100110000111",
		b"111111000110100001111000",
		b"111111001000011111010010",
		b"111111001010011110010001",
		b"111111001100011110101111",
		b"111111001110100000101000",
		b"111111010000100011110110",
		b"111111010010101000010110",
		b"111111010100101110000001",
		b"111111010110110100110011",
		b"111111011000111100100111",
		b"111111011011000101010111",
		b"111111011101001110111111",
		b"111111011111011001011010",
		b"111111100001100100100010",
		b"111111100011110000010010",
		b"111111100101111100100110",
		b"111111101000001001010111",
		b"111111101010010110100010",
		b"111111101100100100000000",
		b"111111101110110001101110",
		b"111111110000111111100101",
		b"111111110011001101100000",
		b"111111110101011011011011",
		b"111111110111101001010000",
		b"111111111001110110111011",
		b"111111111100000100010110",
		b"111111111110010001011101",
		b"000000000000011110001001",
		b"000000000010101010011000",
		b"000000000100110110000011",
		b"000000000111000001000101",
		b"000000001001001011011011",
		b"000000001011010100111111",
		b"000000001101011101101100",
		b"000000001111100101011101",
		b"000000010001101100001111",
		b"000000010011110001111100",
		b"000000010101110110100000",
		b"000000010111111001110111",
		b"000000011001111011111011",
		b"000000011011111100101001",
		b"000000011101111011111101",
		b"000000011111111001110001",
		b"000000100001110110000010",
		b"000000100011110000101100",
		b"000000100101101001101011",
		b"000000100111100000111010",
		b"000000101001010110010110",
		b"000000101011001001111100",
		b"000000101100111011100110",
		b"000000101110101011010011",
		b"000000110000011000111101",
		b"000000110010000100100010",
		b"000000110011101101111110",
		b"000000110101010101001110",
		b"000000110110111010001111",
		b"000000111000011100111101",
		b"000000111001111101010101",
		b"000000111011011011010101",
		b"000000111100110110111010",
		b"000000111110010000000000",
		b"000000111111100110100110",
		b"000001000000111010101000",
		b"000001000010001100000101",
		b"000001000011011010111001",
		b"000001000100100111000010",
		b"000001000101110000011111",
		b"000001000110110111001110",
		b"000001000111111011001011",
		b"000001001000111100010110",
		b"000001001001111010101101",
		b"000001001010110110001101",
		b"000001001011101110110111",
		b"000001001100100100100111",
		b"000001001101010111011101",
		b"000001001110000111010111",
		b"000001001110110100010101",
		b"000001001111011110010101",
		b"000001010000000101010111",
		b"000001010000101001011010",
		b"000001010001001010011100",
		b"000001010001101000011110",
		b"000001010010000011011111",
		b"000001010010011011011111",
		b"000001010010110000011101",
		b"000001010011000010011001",
		b"000001010011010001010100",
		b"000001010011011101001100",
		b"000001010011100110000100",
		b"000001010011101011111010",
		b"000001010011101110101111",
		b"000001010011101110100100",
		b"000001010011101011011010",
		b"000001010011100101010000",
		b"000001010011011100001001",
		b"000001010011010000000100",
		b"000001010011000001000011",
		b"000001010010101111000111",
		b"000001010010011010010001",
		b"000001010010000010100011",
		b"000001010001100111111101",
		b"000001010001001010100010",
		b"000001010000101010010011",
		b"000001010000000111010010",
		b"000001001111100001100001",
		b"000001001110111001000000",
		b"000001001110001101110100",
		b"000001001101011111111101",
		b"000001001100101111011110",
		b"000001001011111100011000",
		b"000001001011000110101111",
		b"000001001010001110100101",
		b"000001001001010011111100",
		b"000001001000010110110111",
		b"000001000111010111011000",
		b"000001000110010101100011",
		b"000001000101010001011010",
		b"000001000100001011000000",
		b"000001000011000010010111",
		b"000001000001110111100100",
		b"000001000000101010101000",
		b"000000111111011011101000",
		b"000000111110001010100111",
		b"000000111100110111100111",
		b"000000111011100010101100",
		b"000000111010001011111010",
		b"000000111000110011010100",
		b"000000110111011000111101",
		b"000000110101111100111001",
		b"000000110100011111001100",
		b"000000110010111111111001",
		b"000000110001011111000101",
		b"000000101111111100110010",
		b"000000101110011001000101",
		b"000000101100110100000001",
		b"000000101011001101101011",
		b"000000101001100110000110",
		b"000000100111111101010110",
		b"000000100110010011011111",
		b"000000100100101000100110",
		b"000000100010111100101101",
		b"000000100001001111111010",
		b"000000011111100010010000",
		b"000000011101110011110011",
		b"000000011100000100101000",
		b"000000011010010100110011",
		b"000000011000100100010111",
		b"000000010110110011011001",
		b"000000010101000001111100",
		b"000000010011010000000110",
		b"000000010001011101111010",
		b"000000001111101011011101",
		b"000000001101111000110010",
		b"000000001100000101111101",
		b"000000001010010011000100",
		b"000000001000100000001001",
		b"000000000110101101010001",
		b"000000000100111010100000",
		b"000000000011000111111011",
		b"000000000001010101100100",
		b"111111111111100011100001",
		b"111111111101110001110101",
		b"111111111100000000100100",
		b"111111111010001111110010",
		b"111111111000011111100100",
		b"111111110110101111111100",
		b"111111110101000001000000",
		b"111111110011010010110010",
		b"111111110001100101010110",
		b"111111101111111000110001",
		b"111111101110001101000110",
		b"111111101100100010011000",
		b"111111101010111000101011",
		b"111111101001010000000100",
		b"111111100111101000100100",
		b"111111100110000010010001",
		b"111111100100011101001100",
		b"111111100010111001011010",
		b"111111100001010110111110",
		b"111111011111110101111100",
		b"111111011110010110010101",
		b"111111011100111000001110",
		b"111111011011011011101010",
		b"111111011010000000101011",
		b"111111011000100111010100",
		b"111111010111001111101001",
		b"111111010101111001101100",
		b"111111010100100101100000",
		b"111111010011010011000111",
		b"111111010010000010100101",
		b"111111010000110011111011",
		b"111111001111100111001100",
		b"111111001110011100011011",
		b"111111001101010011101010",
		b"111111001100001100111010",
		b"111111001011001000001111",
		b"111111001010000101101001",
		b"111111001001000101001100",
		b"111111001000000110111001",
		b"111111000111001010110010",
		b"111111000110010000111000",
		b"111111000101011001001101",
		b"111111000100100011110011",
		b"111111000011110000101100",
		b"111111000010111111111000",
		b"111111000010010001011001",
		b"111111000001100101010000",
		b"111111000000111011011110",
		b"111111000000010100000100",
		b"111110111111101111000100",
		b"111110111111001100011101",
		b"111110111110101100010010",
		b"111110111110001110100010",
		b"111110111101110011001110",
		b"111110111101011010010111",
		b"111110111101000011111101",
		b"111110111100110000000001",
		b"111110111100011110100010",
		b"111110111100001111100000",
		b"111110111100000010111101",
		b"111110111011111000110111",
		b"111110111011110001010000",
		b"111110111011101100000101",
		b"111110111011101001011000",
		b"111110111011101001001000",
		b"111110111011101011010100",
		b"111110111011101111111100",
		b"111110111011110110111111",
		b"111110111100000000011101",
		b"111110111100001100010101",
		b"111110111100011010100101",
		b"111110111100101011001101",
		b"111110111100111110001100",
		b"111110111101010011100001",
		b"111110111101101011001010",
		b"111110111110000101000111",
		b"111110111110100001010101",
		b"111110111110111111110100",
		b"111110111111100000100001",
		b"111111000000000011011100",
		b"111111000000101000100011",
		b"111111000001001111110011",
		b"111111000001111001001100",
		b"111111000010100100101011",
		b"111111000011010010001110",
		b"111111000100000001110011",
		b"111111000100110011011000",
		b"111111000101100110111100",
		b"111111000110011100011011",
		b"111111000111010011110100",
		b"111111001000001101000100",
		b"111111001001001000001001",
		b"111111001010000101000000",
		b"111111001011000011101000",
		b"111111001100000011111100",
		b"111111001101000101111011",
		b"111111001110001001100010",
		b"111111001111001110101110",
		b"111111010000010101011101",
		b"111111010001011101101100",
		b"111111010010100111010111",
		b"111111010011110010011100",
		b"111111010100111110111001",
		b"111111010110001100101001",
		b"111111010111011011101010",
		b"111111011000101011111001",
		b"111111011001111101010100",
		b"111111011011001111110101",
		b"111111011100100011011100",
		b"111111011101111000000011",
		b"111111011111001101101001",
		b"111111100000100100001010",
		b"111111100001111011100011",
		b"111111100011010011110000",
		b"111111100100101100101110",
		b"111111100110000110011010",
		b"111111100111100000110000",
		b"111111101000111011101101",
		b"111111101010010111001110",
		b"111111101011110011010000",
		b"111111101101001111101110",
		b"111111101110101100100110",
		b"111111110000001001110101",
		b"111111110001100111010110",
		b"111111110011000101000110",
		b"111111110100100011000011",
		b"111111110110000001001000",
		b"111111110111011111010011",
		b"111111111000111101011111",
		b"111111111010011011101010",
		b"111111111011111001110000",
		b"111111111101010111101110",
		b"111111111110110101100001",
		b"000000000000010011000100",
		b"000000000001110000010110",
		b"000000000011001101010010",
		b"000000000100101001110110",
		b"000000000110000101111110",
		b"000000000111100001100110",
		b"000000001000111100101101",
		b"000000001010010111001110",
		b"000000001011110001000111",
		b"000000001101001010010100",
		b"000000001110100010110010",
		b"000000001111111010011111",
		b"000000010001010001010111",
		b"000000010010100111010111",
		b"000000010011111100011101",
		b"000000010101010000100110",
		b"000000010110100011101110",
		b"000000010111110101110100",
		b"000000011001000110110100",
		b"000000011010010110101011",
		b"000000011011100101010111",
		b"000000011100110010110110",
		b"000000011101111111000101",
		b"000000011111001010000001",
		b"000000100000010011101000",
		b"000000100001011011110111",
		b"000000100010100010101101",
		b"000000100011101000000110",
		b"000000100100101100000010",
		b"000000100101101110011101",
		b"000000100110101111010101",
		b"000000100111101110101001",
		b"000000101000101100010111",
		b"000000101001101000011100",
		b"000000101010100010110111",
		b"000000101011011011100110",
		b"000000101100010010100111",
		b"000000101101000111111001",
		b"000000101101111011011010",
		b"000000101110101101001000",
		b"000000101111011101000011",
		b"000000110000001011001000",
		b"000000110000110111010111",
		b"000000110001100001101101",
		b"000000110010001010001011",
		b"000000110010110000101111",
		b"000000110011010101011000",
		b"000000110011111000000101",
		b"000000110100011000110101",
		b"000000110100110111100111",
		b"000000110101010100011010",
		b"000000110101101111001111",
		b"000000110110001000000100",
		b"000000110110011110111000",
		b"000000110110110011101100",
		b"000000110111000110011111",
		b"000000110111010111010001",
		b"000000110111100110000001",
		b"000000110111110010101111",
		b"000000110111111101011011",
		b"000000111000000110000110",
		b"000000111000001100101111",
		b"000000111000010001010110",
		b"000000111000010011111100",
		b"000000111000010100100001",
		b"000000111000010011000101",
		b"000000111000001111101001",
		b"000000111000001010001100",
		b"000000111000000010110001",
		b"000000110111111001010111",
		b"000000110111101101111111",
		b"000000110111100000101001",
		b"000000110111010001011000",
		b"000000110111000000001011",
		b"000000110110101101000011",
		b"000000110110011000000010",
		b"000000110110000001001001",
		b"000000110101101000011000",
		b"000000110101001101110001",
		b"000000110100110001010110",
		b"000000110100010011001000",
		b"000000110011110011000111",
		b"000000110011010001010110",
		b"000000110010101101110110",
		b"000000110010001000101001",
		b"000000110001100001110000",
		b"000000110000111001001101",
		b"000000110000001111000010",
		b"000000101111100011010000",
		b"000000101110110101111010",
		b"000000101110000111000001",
		b"000000101101010110100111",
		b"000000101100100100101110",
		b"000000101011110001011001",
		b"000000101010111100101010",
		b"000000101010000110100001",
		b"000000101001001111000011",
		b"000000101000010110010000",
		b"000000100111011100001100",
		b"000000100110100000111000",
		b"000000100101100100010111",
		b"000000100100100110101011",
		b"000000100011100111110111",
		b"000000100010100111111101",
		b"000000100001100111000000",
		b"000000100000100101000001",
		b"000000011111100010000101",
		b"000000011110011110001100",
		b"000000011101011001011011",
		b"000000011100010011110010",
		b"000000011011001101010110",
		b"000000011010000110001000",
		b"000000011000111110001100",
		b"000000010111110101100100",
		b"000000010110101100010010",
		b"000000010101100010011011",
		b"000000010100010111111111",
		b"000000010011001101000010",
		b"000000010010000001101000",
		b"000000010000110101110001",
		b"000000001111101001100010",
		b"000000001110011100111110",
		b"000000001101010000000110",
		b"000000001100000010111110",
		b"000000001010110101101000",
		b"000000001001101000001000",
		b"000000001000011010011111",
		b"000000000111001100110010",
		b"000000000101111111000010",
		b"000000000100110001010011",
		b"000000000011100011100111",
		b"000000000010010110000001",
		b"000000000001001000100100",
		b"111111111111111011010010",
		b"111111111110101110001110",
		b"111111111101100001011011",
		b"111111111100010100111100",
		b"111111111011001000110011",
		b"111111111001111101000011",
		b"111111111000110001101111",
		b"111111110111100110111000",
		b"111111110110011100100011",
		b"111111110101010010110000",
		b"111111110100001001100100",
		b"111111110011000000111111",
		b"111111110001111001000110",
		b"111111110000110001111010",
		b"111111101111101011011101",
		b"111111101110100101110010",
		b"111111101101100000111100",
		b"111111101100011100111101",
		b"111111101011011001110110",
		b"111111101010010111101010",
		b"111111101001010110011100",
		b"111111101000010110001101",
		b"111111100111010111000000",
		b"111111100110011000110111",
		b"111111100101011011110011",
		b"111111100100011111110111",
		b"111111100011100101000101",
		b"111111100010101011011110",
		b"111111100001110011000100",
		b"111111100000111011111010",
		b"111111100000000110000000",
		b"111111011111010001011001",
		b"111111011110011110000110",
		b"111111011101101100001001",
		b"111111011100111011100011",
		b"111111011100001100010110",
		b"111111011011011110100011",
		b"111111011010110010001100",
		b"111111011010000111010010",
		b"111111011001011101110110",
		b"111111011000110101111001",
		b"111111011000001111011101",
		b"111111010111101010100011",
		b"111111010111000111001011",
		b"111111010110100101010111",
		b"111111010110000101000111",
		b"111111010101100110011101",
		b"111111010101001001011010",
		b"111111010100101101111101",
		b"111111010100010100001000",
		b"111111010011111011111011",
		b"111111010011100101011000",
		b"111111010011010000011101",
		b"111111010010111101001101",
		b"111111010010101011100110",
		b"111111010010011011101011",
		b"111111010010001101011010",
		b"111111010010000000110100",
		b"111111010001110101111001",
		b"111111010001101100101010",
		b"111111010001100101000101",
		b"111111010001011111001100",
		b"111111010001011010111111",
		b"111111010001011000011100",
		b"111111010001010111100100",
		b"111111010001011000010111",
		b"111111010001011010110011",
		b"111111010001011110111010",
		b"111111010001100100101010",
		b"111111010001101100000011",
		b"111111010001110101000100",
		b"111111010001111111101101",
		b"111111010010001011111100",
		b"111111010010011001110011",
		b"111111010010101001001110",
		b"111111010010111010001110",
		b"111111010011001100110010",
		b"111111010011100000111001",
		b"111111010011110110100010",
		b"111111010100001101101100",
		b"111111010100100110010101",
		b"111111010101000000011100",
		b"111111010101011100000010",
		b"111111010101111001000011",
		b"111111010110010111011111",
		b"111111010110110111010100",
		b"111111010111011000100010",
		b"111111010111111011000110",
		b"111111011000011110111111",
		b"111111011001000100001100",
		b"111111011001101010101011",
		b"111111011010010010011011",
		b"111111011010111011011001",
		b"111111011011100101100101",
		b"111111011100010000111100",
		b"111111011100111101011101",
		b"111111011101101011000101",
		b"111111011110011001110100",
		b"111111011111001001100111",
		b"111111011111111010011100",
		b"111111100000101100010001",
		b"111111100001011111000101",
		b"111111100010010010110110",
		b"111111100011000111100000",
		b"111111100011111101000100",
		b"111111100100110011011101",
		b"111111100101101010101011",
		b"111111100110100010101011",
		b"111111100111011011011011",
		b"111111101000010100111000",
		b"111111101001001111000001",
		b"111111101010001001110100",
		b"111111101011000101001110",
		b"111111101100000001001101",
		b"111111101100111101101111",
		b"111111101101111010110001",
		b"111111101110111000010010",
		b"111111101111110110001110",
		b"111111110000110100100100",
		b"111111110001110011010010",
		b"111111110010110010010101",
		b"111111110011110001101010",
		b"111111110100110001010000",
		b"111111110101110001000100",
		b"111111110110110001000100",
		b"111111110111110001001110",
		b"111111111000110001011110",
		b"111111111001110001110100",
		b"111111111010110010001100",
		b"111111111011110010100101",
		b"111111111100110010111100",
		b"111111111101110011001110",
		b"111111111110110011011010",
		b"111111111111110011011101",
		b"000000000000110011010101",
		b"000000000001110011000000",
		b"000000000010110010011011",
		b"000000000011110001100101",
		b"000000000100110000011010",
		b"000000000101101110111010",
		b"000000000110101101000001",
		b"000000000111101010101101",
		b"000000001000100111111101",
		b"000000001001100100101111",
		b"000000001010100001000000",
		b"000000001011011100101110",
		b"000000001100010111110111",
		b"000000001101010010011001",
		b"000000001110001100010011",
		b"000000001111000101100010",
		b"000000001111111110000100",
		b"000000010000110101111000",
		b"000000010001101100111011",
		b"000000010010100011001100",
		b"000000010011011000101001",
		b"000000010100001101010000",
		b"000000010101000001000000",
		b"000000010101110011110111",
		b"000000010110100101110010",
		b"000000010111010110110010",
		b"000000011000000110110011",
		b"000000011000110101110101",
		b"000000011001100011110110",
		b"000000011010010000110100",
		b"000000011010111100101111",
		b"000000011011100111100100",
		b"000000011100010001010010",
		b"000000011100111001111001",
		b"000000011101100001010110",
		b"000000011110000111101010",
		b"000000011110101100110001",
		b"000000011111010000101100",
		b"000000011111110011011010",
		b"000000100000010100111001",
		b"000000100000110101001000",
		b"000000100001010100000110",
		b"000000100001110001110100",
		b"000000100010001110001110",
		b"000000100010101001010110",
		b"000000100011000011001010",
		b"000000100011011011101010",
		b"000000100011110010110100",
		b"000000100100001000101001",
		b"000000100100011101001000",
		b"000000100100110000010000",
		b"000000100101000010000000",
		b"000000100101010010011001",
		b"000000100101100001011011",
		b"000000100101101111000100",
		b"000000100101111011010101",
		b"000000100110000110001101",
		b"000000100110001111101101",
		b"000000100110010111110011",
		b"000000100110011110100001",
		b"000000100110100011110110",
		b"000000100110100111110011",
		b"000000100110101010010110",
		b"000000100110101011100001",
		b"000000100110101011010100",
		b"000000100110101001101111",
		b"000000100110100110110010",
		b"000000100110100010011110",
		b"000000100110011100110011",
		b"000000100110010101110001",
		b"000000100110001101011001",
		b"000000100110000011101100",
		b"000000100101111000101010",
		b"000000100101101100010011",
		b"000000100101011110101001",
		b"000000100101001111101100",
		b"000000100100111111011101",
		b"000000100100101101111100",
		b"000000100100011011001100",
		b"000000100100000111001011",
		b"000000100011110001111100",
		b"000000100011011011100000",
		b"000000100011000011110110",
		b"000000100010101011000001",
		b"000000100010010001000010",
		b"000000100001110101111001",
		b"000000100001011001101001",
		b"000000100000111100010001",
		b"000000100000011101110011",
		b"000000011111111110010001",
		b"000000011111011101101100",
		b"000000011110111100000101",
		b"000000011110011001011110",
		b"000000011101110101111000",
		b"000000011101010001010100",
		b"000000011100101011110101",
		b"000000011100000101011010",
		b"000000011011011110000111",
		b"000000011010110101111100",
		b"000000011010001100111011",
		b"000000011001100011000110",
		b"000000011000111000011111",
		b"000000011000001101000110",
		b"000000010111100000111110",
		b"000000010110110100001001",
		b"000000010110000110100111",
		b"000000010101011000011100",
		b"000000010100101001101000",
		b"000000010011111010001110",
		b"000000010011001010001111",
		b"000000010010011001101100",
		b"000000010001101000101001",
		b"000000010000110111000110",
		b"000000010000000101000110",
		b"000000001111010010101011",
		b"000000001110011111110101",
		b"000000001101101100101000",
		b"000000001100111001000101",
		b"000000001100000101001101",
		b"000000001011010001000100",
		b"000000001010011100101010",
		b"000000001001101000000010",
		b"000000001000110011001101",
		b"000000000111111110001110",
		b"000000000111001001000110",
		b"000000000110010011111000",
		b"000000000101011110100101",
		b"000000000100101001001111",
		b"000000000011110011110111",
		b"000000000010111110100001",
		b"000000000010001001001110",
		b"000000000001010011111111",
		b"000000000000011110110111",
		b"111111111111101001111000",
		b"111111111110110101000010",
		b"111111111110000000011001",
		b"111111111101001011111110",
		b"111111111100010111110011",
		b"111111111011100011111001",
		b"111111111010110000010011",
		b"111111111001111101000010",
		b"111111111001001010001000",
		b"111111111000010111100110",
		b"111111110111100101100000",
		b"111111110110110011110101",
		b"111111110110000010101000",
		b"111111110101010001111011",
		b"111111110100100001101110",
		b"111111110011110010000101",
		b"111111110011000011000000",
		b"111111110010010100100000",
		b"111111110001100110101001",
		b"111111110000111001011010",
		b"111111110000001100110110",
		b"111111101111100000111101",
		b"111111101110110101110010",
		b"111111101110001011010110",
		b"111111101101100001101010",
		b"111111101100111000110000",
		b"111111101100010000101000",
		b"111111101011101001010100",
		b"111111101011000010110110",
		b"111111101010011101001111",
		b"111111101001111000011111",
		b"111111101001010100101000",
		b"111111101000110001101011",
		b"111111101000001111101001",
		b"111111100111101110100011",
		b"111111100111001110011011",
		b"111111100110101111010000",
		b"111111100110010001000101",
		b"111111100101110011111001",
		b"111111100101010111101110",
		b"111111100100111100100101",
		b"111111100100100010011111",
		b"111111100100001001011011",
		b"111111100011110001011011",
		b"111111100011011010100000",
		b"111111100011000100101010",
		b"111111100010101111111001",
		b"111111100010011100001111",
		b"111111100010001001101100",
		b"111111100001111000001111",
		b"111111100001100111111011",
		b"111111100001011000101110",
		b"111111100001001010101001",
		b"111111100000111101101110",
		b"111111100000110001111011",
		b"111111100000100111010001",
		b"111111100000011101110000",
		b"111111100000010101011001",
		b"111111100000001110001011",
		b"111111100000001000000111",
		b"111111100000000011001100",
		b"111111011111111111011011",
		b"111111011111111100110011",
		b"111111011111111011010101",
		b"111111011111111010111111",
		b"111111011111111011110011",
		b"111111011111111101101111",
		b"111111100000000000110100",
		b"111111100000000101000001",
		b"111111100000001010010101",
		b"111111100000010000110001",
		b"111111100000011000010100",
		b"111111100000100000111110",
		b"111111100000101010101101",
		b"111111100000110101100010",
		b"111111100001000001011100",
		b"111111100001001110011010",
		b"111111100001011100011011",
		b"111111100001101011011111",
		b"111111100001111011100110",
		b"111111100010001100101110",
		b"111111100010011110110110",
		b"111111100010110001111111",
		b"111111100011000110000110",
		b"111111100011011011001011",
		b"111111100011110001001101",
		b"111111100100001000001100",
		b"111111100100100000000101",
		b"111111100100111000111001",
		b"111111100101010010100110",
		b"111111100101101101001011",
		b"111111100110001000100110",
		b"111111100110100100111000",
		b"111111100111000001111110",
		b"111111100111011111111000",
		b"111111100111111110100100",
		b"111111101000011110000000",
		b"111111101000111110001101",
		b"111111101001011111001000",
		b"111111101010000000110000",
		b"111111101010100011000100",
		b"111111101011000110000011",
		b"111111101011101001101010",
		b"111111101100001101111010",
		b"111111101100110010110000",
		b"111111101101011000001010",
		b"111111101101111110001001",
		b"111111101110100100101001",
		b"111111101111001011101010",
		b"111111101111110011001010",
		b"111111110000011011000111",
		b"111111110001000011100001",
		b"111111110001101100010101",
		b"111111110010010101100011",
		b"111111110010111111001000",
		b"111111110011101001000011",
		b"111111110100010011010010",
		b"111111110100111101110101",
		b"111111110101101000101000",
		b"111111110110010011101100",
		b"111111110110111110111101",
		b"111111110111101010011011",
		b"111111111000010110000101",
		b"111111111001000001110111",
		b"111111111001101101110010",
		b"111111111010011001110011",
		b"111111111011000101111000",
		b"111111111011110010000001",
		b"111111111100011110001011",
		b"111111111101001010010110",
		b"111111111101110110011110",
		b"111111111110100010100100",
		b"111111111111001110100101",
		b"111111111111111010011111",
		b"000000000000100110010010",
		b"000000000001010001111100",
		b"000000000001111101011010",
		b"000000000010101000101100",
		b"000000000011010011110001",
		b"000000000011111110100110",
		b"000000000100101001001010",
		b"000000000101010011011100",
		b"000000000101111101011011",
		b"000000000110100111000100",
		b"000000000111010000010110",
		b"000000000111111001010001",
		b"000000001000100001110010",
		b"000000001001001001111000",
		b"000000001001110001100011",
		b"000000001010011000110000",
		b"000000001010111111011110",
		b"000000001011100101101101",
		b"000000001100001011011010",
		b"000000001100110000100100",
		b"000000001101010101001011",
		b"000000001101111001001101",
		b"000000001110011100101001",
		b"000000001110111111011101",
		b"000000001111100001101010",
		b"000000010000000011001100",
		b"000000010000100100000101",
		b"000000010001000100010010",
		b"000000010001100011110010",
		b"000000010010000010100100",
		b"000000010010100000101000",
		b"000000010010111101111101",
		b"000000010011011010100001",
		b"000000010011110110010100",
		b"000000010100010001010101",
		b"000000010100101011100011",
		b"000000010101000100111101",
		b"000000010101011101100011",
		b"000000010101110101010100",
		b"000000010110001100001110",
		b"000000010110100010010011",
		b"000000010110110111100000",
		b"000000010111001011110101",
		b"000000010111011111010010",
		b"000000010111110001110111",
		b"000000011000000011100010",
		b"000000011000010100010011",
		b"000000011000100100001010",
		b"000000011000110011000110",
		b"000000011001000001001000",
		b"000000011001001110001110",
		b"000000011001011010011001",
		b"000000011001100101100111",
		b"000000011001101111111010",
		b"000000011001111001010000",
		b"000000011010000001101010",
		b"000000011010001001001000",
		b"000000011010001111101001",
		b"000000011010010101001101",
		b"000000011010011001110100",
		b"000000011010011101011111",
		b"000000011010100000001101",
		b"000000011010100001111110",
		b"000000011010100010110100",
		b"000000011010100010101100",
		b"000000011010100001101001",
		b"000000011010011111101001",
		b"000000011010011100101110",
		b"000000011010011000111000",
		b"000000011010010100000110",
		b"000000011010001110011010",
		b"000000011010000111110011",
		b"000000011010000000010010",
		b"000000011001110111111000",
		b"000000011001101110100101",
		b"000000011001100100011001",
		b"000000011001011001010101",
		b"000000011001001101011001",
		b"000000011001000000100111",
		b"000000011000110010111110",
		b"000000011000100100011111",
		b"000000011000010101001100",
		b"000000011000000101000100",
		b"000000010111110100001000",
		b"000000010111100010011010",
		b"000000010111001111111010",
		b"000000010110111100101000",
		b"000000010110101000100110",
		b"000000010110010011110100",
		b"000000010101111110010011",
		b"000000010101101000000101",
		b"000000010101010001001010",
		b"000000010100111001100011",
		b"000000010100100001010001",
		b"000000010100001000010100",
		b"000000010011101110101111",
		b"000000010011010100100010",
		b"000000010010111001101110",
		b"000000010010011110010100",
		b"000000010010000010010101",
		b"000000010001100101110011",
		b"000000010001001000101101",
		b"000000010000101011000111",
		b"000000010000001101000000",
		b"000000001111101110011010",
		b"000000001111001111010110",
		b"000000001110101111110101",
		b"000000001110001111111001",
		b"000000001101101111100010",
		b"000000001101001110110010",
		b"000000001100101101101010",
		b"000000001100001100001100",
		b"000000001011101010011000",
		b"000000001011001000001111",
		b"000000001010100101110100",
		b"000000001010000011001000",
		b"000000001001100000001011",
		b"000000001000111100111110",
		b"000000001000011001100101",
		b"000000000111110101111110",
		b"000000000111010010001101",
		b"000000000110101110010001",
		b"000000000110001010001101",
		b"000000000101100110000010",
		b"000000000101000001110001",
		b"000000000100011101011011",
		b"000000000011111001000001",
		b"000000000011010100100110",
		b"000000000010110000001010",
		b"000000000010001011101110",
		b"000000000001100111010100",
		b"000000000001000010111101",
		b"000000000000011110101011",
		b"111111111111111010011110",
		b"111111111111010110011000",
		b"111111111110110010011010",
		b"111111111110001110100110",
		b"111111111101101010111100",
		b"111111111101000111011110",
		b"111111111100100100001110",
		b"111111111100000001001011",
		b"111111111011011110011000",
		b"111111111010111011110110",
		b"111111111010011001100110",
		b"111111111001110111101000",
		b"111111111001010101111111",
		b"111111111000110100101011",
		b"111111111000010011101110",
		b"111111110111110011001000",
		b"111111110111010010111010",
		b"111111110110110011000111",
		b"111111110110010011101110",
		b"111111110101110100110000",
		b"111111110101010110010000",
		b"111111110100111000001101",
		b"111111110100011010101001",
		b"111111110011111101100101",
		b"111111110011100001000010",
		b"111111110011000101000000",
		b"111111110010101001100000",
		b"111111110010001110100100",
		b"111111110001110100001100",
		b"111111110001011010011001",
		b"111111110001000001001011",
		b"111111110000101000100101",
		b"111111110000010000100101",
		b"111111101111111001001110",
		b"111111101111100010011111",
		b"111111101111001100011010",
		b"111111101110110110111111",
		b"111111101110100010001111",
		b"111111101110001110001010",
		b"111111101101111010110001",
		b"111111101101101000000101",
		b"111111101101010110000110",
		b"111111101101000100110100",
		b"111111101100110100010000",
		b"111111101100100100011011",
		b"111111101100010101010101",
		b"111111101100000110111110",
		b"111111101011111001010110",
		b"111111101011101100011111",
		b"111111101011100000011000",
		b"111111101011010101000001",
		b"111111101011001010011011",
		b"111111101011000000100111",
		b"111111101010110111100100",
		b"111111101010101111010010",
		b"111111101010100111110010",
		b"111111101010100001000011",
		b"111111101010011011000111",
		b"111111101010010101111100",
		b"111111101010010001100011",
		b"111111101010001101111100",
		b"111111101010001011000111",
		b"111111101010001001000100",
		b"111111101010000111110011",
		b"111111101010000111010011",
		b"111111101010000111100101",
		b"111111101010001000101001",
		b"111111101010001010011101",
		b"111111101010001101000011",
		b"111111101010010000011010",
		b"111111101010010100100000",
		b"111111101010011001011000",
		b"111111101010011110111111",
		b"111111101010100101010101",
		b"111111101010101100011011",
		b"111111101010110100010000",
		b"111111101010111100110011",
		b"111111101011000110000100",
		b"111111101011010000000011",
		b"111111101011011010101111",
		b"111111101011100110000111",
		b"111111101011110010001011",
		b"111111101011111110111010",
		b"111111101100001100010101",
		b"111111101100011010011001",
		b"111111101100101001000111",
		b"111111101100111000011111",
		b"111111101101001000011110",
		b"111111101101011001000101",
		b"111111101101101010010011",
		b"111111101101111100001000",
		b"111111101110001110100001",
		b"111111101110100001100000",
		b"111111101110110101000010",
		b"111111101111001001000111",
		b"111111101111011101101111",
		b"111111101111110010111000",
		b"111111110000001000100010",
		b"111111110000011110101100",
		b"111111110000110101010100",
		b"111111110001001100011011",
		b"111111110001100011111110",
		b"111111110001111011111110",
		b"111111110010010100011001",
		b"111111110010101101001110",
		b"111111110011000110011101",
		b"111111110011100000000100",
		b"111111110011111010000010",
		b"111111110100010100010111",
		b"111111110100101111000010",
		b"111111110101001010000000",
		b"111111110101100101010010",
		b"111111110110000000110111",
		b"111111110110011100101101",
		b"111111110110111000110011",
		b"111111110111010101001000",
		b"111111110111110001101100",
		b"111111111000001110011100",
		b"111111111000101011011001",
		b"111111111001001000100001",
		b"111111111001100101110011",
		b"111111111010000011001110",
		b"111111111010100000110001",
		b"111111111010111110011010",
		b"111111111011011100001010",
		b"111111111011111001111110",
		b"111111111100010111110101",
		b"111111111100110101101111",
		b"111111111101010011101011",
		b"111111111101110001100111",
		b"111111111110001111100010",
		b"111111111110101101011100",
		b"111111111111001011010011",
		b"111111111111101001000110",
		b"000000000000000110110100",
		b"000000000000100100011101",
		b"000000000001000001111110",
		b"000000000001011111011000",
		b"000000000001111100101000",
		b"000000000010011001101111",
		b"000000000010110110101011",
		b"000000000011010011011011",
		b"000000000011101111111110",
		b"000000000100001100010011",
		b"000000000100101000011001",
		b"000000000101000100001111",
		b"000000000101011111110101",
		b"000000000101111011001001",
		b"000000000110010110001011",
		b"000000000110110000111001",
		b"000000000111001011010010",
		b"000000000111100101010111",
		b"000000000111111111000101",
		b"000000001000011000011101",
		b"000000001000110001011101",
		b"000000001001001010000100",
		b"000000001001100010010010",
		b"000000001001111010000110",
		b"000000001010010001011111",
		b"000000001010101000011100",
		b"000000001010111110111101",
		b"000000001011010101000001",
		b"000000001011101010100111",
		b"000000001011111111101111",
		b"000000001100010100010111",
		b"000000001100101000100000",
		b"000000001100111100001001",
		b"000000001101001111010000",
		b"000000001101100001110111",
		b"000000001101110011111011",
		b"000000001110000101011100",
		b"000000001110010110011011",
		b"000000001110100110110101",
		b"000000001110110110101100",
		b"000000001111000101111110",
		b"000000001111010100101100",
		b"000000001111100010110100",
		b"000000001111110000010110",
		b"000000001111111101010010",
		b"000000010000001001101000",
		b"000000010000010101010110",
		b"000000010000100000011110",
		b"000000010000101010111111",
		b"000000010000110100111000",
		b"000000010000111110001001",
		b"000000010001000110110010",
		b"000000010001001110110010",
		b"000000010001010110001011",
		b"000000010001011100111011",
		b"000000010001100011000010",
		b"000000010001101000100001",
		b"000000010001101101010110",
		b"000000010001110001100011",
		b"000000010001110101000111",
		b"000000010001111000000011",
		b"000000010001111010010101",
		b"000000010001111011111111",
		b"000000010001111100111111",
		b"000000010001111101011000",
		b"000000010001111101000111",
		b"000000010001111100001111",
		b"000000010001111010101101",
		b"000000010001111000100100",
		b"000000010001110101110011",
		b"000000010001110010011011",
		b"000000010001101110011011",
		b"000000010001101001110011",
		b"000000010001100100100101",
		b"000000010001011110110001",
		b"000000010001011000010110",
		b"000000010001010001010101",
		b"000000010001001001101110",
		b"000000010001000001100011",
		b"000000010000111000110010",
		b"000000010000101111011110",
		b"000000010000100101100101",
		b"000000010000011011001001",
		b"000000010000010000001010",
		b"000000010000000100101000",
		b"000000001111111000100101",
		b"000000001111101100000000",
		b"000000001111011110111010",
		b"000000001111010001010100",
		b"000000001111000011001110",
		b"000000001110110100101000",
		b"000000001110100101100101",
		b"000000001110010110000011",
		b"000000001110000110000100",
		b"000000001101110101101000",
		b"000000001101100100110001",
		b"000000001101010011011110",
		b"000000001101000001110000",
		b"000000001100101111101001",
		b"000000001100011101001000",
		b"000000001100001010001111",
		b"000000001011110110111110",
		b"000000001011100011010111",
		b"000000001011001111011001",
		b"000000001010111011000101",
		b"000000001010100110011101",
		b"000000001010010001100001",
		b"000000001001111100010010",
		b"000000001001100110110001",
		b"000000001001010000111110",
		b"000000001000111010111011",
		b"000000001000100100100111",
		b"000000001000001110000101",
		b"000000000111110111010101",
		b"000000000111100000010111",
		b"000000000111001001001101",
		b"000000000110110001111000",
		b"000000000110011010010111",
		b"000000000110000010101101",
		b"000000000101101010111010",
		b"000000000101010010111110",
		b"000000000100111010111100",
		b"000000000100100010110011",
		b"000000000100001010100100",
		b"000000000011110010010001",
		b"000000000011011001111010",
		b"000000000011000001100000",
		b"000000000010101001000100",
		b"000000000010010000100111",
		b"000000000001111000001001",
		b"000000000001011111101100",
		b"000000000001000111010001",
		b"000000000000101110110111",
		b"000000000000010110100001",
		b"111111111111111110001111",
		b"111111111111100110000001",
		b"111111111111001101111001",
		b"111111111110110101111000",
		b"111111111110011101111110",
		b"111111111110000110001100",
		b"111111111101101110100011",
		b"111111111101010111000011",
		b"111111111100111111101110",
		b"111111111100101000100101",
		b"111111111100010001100111",
		b"111111111011111010110111",
		b"111111111011100100010011",
		b"111111111011001101111111",
		b"111111111010110111111001",
		b"111111111010100010000100",
		b"111111111010001100011110",
		b"111111111001110111001010",
		b"111111111001100010001000",
		b"111111111001001101011001",
		b"111111111000111000111101",
		b"111111111000100100110101",
		b"111111111000010001000010",
		b"111111110111111101100100",
		b"111111110111101010011011",
		b"111111110111010111101010",
		b"111111110111000101001111",
		b"111111110110110011001100",
		b"111111110110100001100001",
		b"111111110110010000001111",
		b"111111110101111111010110",
		b"111111110101101110110111",
		b"111111110101011110110011",
		b"111111110101001111001001",
		b"111111110100111111111010",
		b"111111110100110001000111",
		b"111111110100100010110000",
		b"111111110100010100110110",
		b"111111110100000111011001",
		b"111111110011111010011001",
		b"111111110011101101110110",
		b"111111110011100001110010",
		b"111111110011010110001100",
		b"111111110011001011000101",
		b"111111110011000000011101",
		b"111111110010110110010100",
		b"111111110010101100101011",
		b"111111110010100011100001",
		b"111111110010011010111000",
		b"111111110010010010101111",
		b"111111110010001011000110",
		b"111111110010000011111101",
		b"111111110001111101010101",
		b"111111110001110111001111",
		b"111111110001110001101001",
		b"111111110001101100100100",
		b"111111110001101000000000",
		b"111111110001100011111101",
		b"111111110001100000011100",
		b"111111110001011101011100",
		b"111111110001011010111101",
		b"111111110001011000111111",
		b"111111110001010111100011",
		b"111111110001010110100111",
		b"111111110001010110001101",
		b"111111110001010110010100",
		b"111111110001010110111011",
		b"111111110001011000000011",
		b"111111110001011001101100",
		b"111111110001011011110110",
		b"111111110001011110011111",
		b"111111110001100001101001",
		b"111111110001100101010010",
		b"111111110001101001011011",
		b"111111110001101110000100",
		b"111111110001110011001011",
		b"111111110001111000110010",
		b"111111110001111110110111",
		b"111111110010000101011010",
		b"111111110010001100011011",
		b"111111110010010011111010",
		b"111111110010011011110110",
		b"111111110010100100001111",
		b"111111110010101101000100",
		b"111111110010110110010110",
		b"111111110011000000000011",
		b"111111110011001010001011",
		b"111111110011010100101110",
		b"111111110011011111101100",
		b"111111110011101011000011",
		b"111111110011110110110100",
		b"111111110100000010111101",
		b"111111110100001111011111",
		b"111111110100011100011001",
		b"111111110100101001101011",
		b"111111110100110111010011",
		b"111111110101000101010001",
		b"111111110101010011100101",
		b"111111110101100010001110",
		b"111111110101110001001100",
		b"111111110110000000011101",
		b"111111110110010000000010",
		b"111111110110011111111010",
		b"111111110110110000000100",
		b"111111110111000000011111",
		b"111111110111010001001100",
		b"111111110111100010001000",
		b"111111110111110011010100",
		b"111111111000000100101111",
		b"111111111000010110011001",
		b"111111111000101000010000",
		b"111111111000111010010100",
		b"111111111001001100100100",
		b"111111111001011111000000",
		b"111111111001110001100110",
		b"111111111010000100010111",
		b"111111111010010111010010",
		b"111111111010101010010101",
		b"111111111010111101100001",
		b"111111111011010000110100",
		b"111111111011100100001101",
		b"111111111011110111101101",
		b"111111111100001011010010",
		b"111111111100011110111100",
		b"111111111100110010101010",
		b"111111111101000110011010",
		b"111111111101011010001110",
		b"111111111101101110000011",
		b"111111111110000001111010",
		b"111111111110010101110000",
		b"111111111110101001100111",
		b"111111111110111101011101",
		b"111111111111010001010001",
		b"111111111111100101000010",
		b"111111111111111000110001",
		b"000000000000001100011100",
		b"000000000000100000000010",
		b"000000000000110011100100",
		b"000000000001000110111111",
		b"000000000001011010010101",
		b"000000000001101101100011",
		b"000000000010000000101001",
		b"000000000010010011101000",
		b"000000000010100110011101",
		b"000000000010111001001000",
		b"000000000011001011101010",
		b"000000000011011110000000",
		b"000000000011110000001011",
		b"000000000100000010001010",
		b"000000000100010011111100",
		b"000000000100100101100010",
		b"000000000100110110111001",
		b"000000000101001000000010",
		b"000000000101011000111100",
		b"000000000101101001100110",
		b"000000000101111010000000",
		b"000000000110001010001010",
		b"000000000110011010000011",
		b"000000000110101001101011",
		b"000000000110111001000000",
		b"000000000111001000000011",
		b"000000000111010110110010",
		b"000000000111100101001111",
		b"000000000111110011010111",
		b"000000001000000001001011",
		b"000000001000001110101010",
		b"000000001000011011110101",
		b"000000001000101000101001",
		b"000000001000110101001000",
		b"000000001001000001010000",
		b"000000001001001101000010",
		b"000000001001011000011101",
		b"000000001001100011100001",
		b"000000001001101110001100",
		b"000000001001111000100000",
		b"000000001010000010011100",
		b"000000001010001100000000",
		b"000000001010010101001010",
		b"000000001010011101111100",
		b"000000001010100110010100",
		b"000000001010101110010011",
		b"000000001010110101111001",
		b"000000001010111101000100",
		b"000000001011000011110110",
		b"000000001011001010001101",
		b"000000001011010000001011",
		b"000000001011010101101110",
		b"000000001011011010110110",
		b"000000001011011111100100",
		b"000000001011100011110111",
		b"000000001011100111101111",
		b"000000001011101011001101",
		b"000000001011101110010000",
		b"000000001011110000111000",
		b"000000001011110011000101",
		b"000000001011110100110111",
		b"000000001011110110001111",
		b"000000001011110111001100",
		b"000000001011110111101110",
		b"000000001011110111110101",
		b"000000001011110111100010",
		b"000000001011110110110101",
		b"000000001011110101101101",
		b"000000001011110100001010",
		b"000000001011110010001110",
		b"000000001011101111111000",
		b"000000001011101101001000",
		b"000000001011101001111110",
		b"000000001011100110011011",
		b"000000001011100010011111",
		b"000000001011011110001010",
		b"000000001011011001011100",
		b"000000001011010100010110",
		b"000000001011001110110111",
		b"000000001011001001000000",
		b"000000001011000010110010",
		b"000000001010111100001100",
		b"000000001010110101001111",
		b"000000001010101101111100",
		b"000000001010100110010010",
		b"000000001010011110010001",
		b"000000001010010101111011",
		b"000000001010001101010000",
		b"000000001010000100010000",
		b"000000001001111010111011",
		b"000000001001110001010010",
		b"000000001001100111010101",
		b"000000001001011101000100",
		b"000000001001010010100001",
		b"000000001001000111101010",
		b"000000001000111100100010",
		b"000000001000110001001000",
		b"000000001000100101011101",
		b"000000001000011001100001",
		b"000000001000001101010101",
		b"000000001000000000111001",
		b"000000000111110100001110",
		b"000000000111100111010011",
		b"000000000111011010001011",
		b"000000000111001100110100",
		b"000000000110111111010001",
		b"000000000110110001100000",
		b"000000000110100011100011",
		b"000000000110010101011011",
		b"000000000110000111000111",
		b"000000000101111000101001",
		b"000000000101101010000000",
		b"000000000101011011001110",
		b"000000000101001100010010",
		b"000000000100111101001110",
		b"000000000100101110000011",
		b"000000000100011110110000",
		b"000000000100001111010101",
		b"000000000011111111110101",
		b"000000000011110000001111",
		b"000000000011100000100100",
		b"000000000011010000110100",
		b"000000000011000001000000",
		b"000000000010110001001001",
		b"000000000010100001001111",
		b"000000000010010001010010",
		b"000000000010000001010100",
		b"000000000001110001010101",
		b"000000000001100001010101",
		b"000000000001010001010100",
		b"000000000001000001010101",
		b"000000000000110001010110",
		b"000000000000100001011001",
		b"000000000000010001011110",
		b"000000000000000001100110",
		b"111111111111110001110001",
		b"111111111111100001111111",
		b"111111111111010010010010",
		b"111111111111000010101010",
		b"111111111110110011000111",
		b"111111111110100011101011",
		b"111111111110010100010100",
		b"111111111110000101000101",
		b"111111111101110101111101",
		b"111111111101100110111101",
		b"111111111101011000000101",
		b"111111111101001001010110",
		b"111111111100111010110001",
		b"111111111100101100010101",
		b"111111111100011110000100",
		b"111111111100001111111110",
		b"111111111100000010000011",
		b"111111111011110100010100",
		b"111111111011100110110001",
		b"111111111011011001011010",
		b"111111111011001100010001",
		b"111111111010111111010101",
		b"111111111010110010100111",
		b"111111111010100110000111",
		b"111111111010011001110110",
		b"111111111010001101110011",
		b"111111111010000010000001",
		b"111111111001110110011110",
		b"111111111001101011001011",
		b"111111111001100000001000",
		b"111111111001010101010110",
		b"111111111001001010110110",
		b"111111111001000000100110",
		b"111111111000110110101001",
		b"111111111000101100111101",
		b"111111111000100011100100",
		b"111111111000011010011101",
		b"111111111000010001101001",
		b"111111111000001001001000",
		b"111111111000000000111010",
		b"111111110111111001000000",
		b"111111110111110001011001",
		b"111111110111101010000110",
		b"111111110111100011001000",
		b"111111110111011100011110",
		b"111111110111010110001000",
		b"111111110111010000000110",
		b"111111110111001010011010",
		b"111111110111000101000010",
		b"111111110110111111111111",
		b"111111110110111011010001",
		b"111111110110110110111001",
		b"111111110110110010110110",
		b"111111110110101111001000",
		b"111111110110101011101111",
		b"111111110110101000101100",
		b"111111110110100101111110",
		b"111111110110100011100110",
		b"111111110110100001100011",
		b"111111110110011111110110",
		b"111111110110011110011110",
		b"111111110110011101011100",
		b"111111110110011100101111",
		b"111111110110011100011000",
		b"111111110110011100010101",
		b"111111110110011100101001",
		b"111111110110011101010001",
		b"111111110110011110001110",
		b"111111110110011111100000",
		b"111111110110100001000111",
		b"111111110110100011000011",
		b"111111110110100101010100",
		b"111111110110100111111001",
		b"111111110110101010110010",
		b"111111110110101101111111",
		b"111111110110110001100000",
		b"111111110110110101010101",
		b"111111110110111001011110",
		b"111111110110111101111010",
		b"111111110111000010101001",
		b"111111110111000111101011",
		b"111111110111001100111111",
		b"111111110111010010100110",
		b"111111110111011000011111",
		b"111111110111011110101010",
		b"111111110111100101000111",
		b"111111110111101011110101",
		b"111111110111110010110100",
		b"111111110111111010000100",
		b"111111111000000001100100",
		b"111111111000001001010100",
		b"111111111000010001010100",
		b"111111111000011001100100",
		b"111111111000100010000010",
		b"111111111000101010110000",
		b"111111111000110011101011",
		b"111111111000111100110101",
		b"111111111001000110001101",
		b"111111111001001111110010",
		b"111111111001011001100100",
		b"111111111001100011100010",
		b"111111111001101101101100",
		b"111111111001111000000011",
		b"111111111010000010100101",
		b"111111111010001101010001",
		b"111111111010011000001000",
		b"111111111010100011001010",
		b"111111111010101110010101",
		b"111111111010111001101010",
		b"111111111011000101000111",
		b"111111111011010000101101",
		b"111111111011011100011011",
		b"111111111011101000010000",
		b"111111111011110100001101",
		b"111111111100000000010000",
		b"111111111100001100011010",
		b"111111111100011000101001",
		b"111111111100100100111110",
		b"111111111100110001011000",
		b"111111111100111101110110",
		b"111111111101001010011000",
		b"111111111101010110111110",
		b"111111111101100011100111",
		b"111111111101110000010011",
		b"111111111101111101000001",
		b"111111111110001001110001",
		b"111111111110010110100010",
		b"111111111110100011010100",
		b"111111111110110000000111",
		b"111111111110111100111001",
		b"111111111111001001101011",
		b"111111111111010110011100",
		b"111111111111100011001100",
		b"111111111111101111111011",
		b"111111111111111100100111",
		b"000000000000001001010000",
		b"000000000000010101110110",
		b"000000000000100010011001",
		b"000000000000101110111000",
		b"000000000000111011010011",
		b"000000000001000111101000",
		b"000000000001010011111001",
		b"000000000001100000000100",
		b"000000000001101100001010",
		b"000000000001111000001000",
		b"000000000010000100000001",
		b"000000000010001111110001",
		b"000000000010011011011011",
		b"000000000010100110111100",
		b"000000000010110010010110",
		b"000000000010111101100110",
		b"000000000011001000101110",
		b"000000000011010011101100",
		b"000000000011011110100000",
		b"000000000011101001001011",
		b"000000000011110011101011",
		b"000000000011111110000000",
		b"000000000100001000001011",
		b"000000000100010010001010",
		b"000000000100011011111101",
		b"000000000100100101100100",
		b"000000000100101110111111",
		b"000000000100111000001110",
		b"000000000101000001001111",
		b"000000000101001010000100",
		b"000000000101010010101011",
		b"000000000101011011000101",
		b"000000000101100011010001",
		b"000000000101101011001111",
		b"000000000101110010111110",
		b"000000000101111010011111",
		b"000000000110000001110001",
		b"000000000110001000110101",
		b"000000000110001111101001",
		b"000000000110010110001101",
		b"000000000110011100100011",
		b"000000000110100010101000",
		b"000000000110101000011110",
		b"000000000110101110000100",
		b"000000000110110011011010",
		b"000000000110111000011111",
		b"000000000110111101010100",
		b"000000000111000001111001",
		b"000000000111000110001101",
		b"000000000111001010010001",
		b"000000000111001110000100",
		b"000000000111010001100101",
		b"000000000111010100110110",
		b"000000000111010111110111",
		b"000000000111011010100110",
		b"000000000111011101000100",
		b"000000000111011111010001",
		b"000000000111100001001101",
		b"000000000111100010111000",
		b"000000000111100100010010",
		b"000000000111100101011010",
		b"000000000111100110010010",
		b"000000000111100110111001",
		b"000000000111100111001110",
		b"000000000111100111010011",
		b"000000000111100111000111",
		b"000000000111100110101010",
		b"000000000111100101111101",
		b"000000000111100100111111",
		b"000000000111100011110000",
		b"000000000111100010010000",
		b"000000000111100000100001",
		b"000000000111011110100001",
		b"000000000111011100010001",
		b"000000000111011001110001",
		b"000000000111010111000001",
		b"000000000111010100000010",
		b"000000000111010000110011",
		b"000000000111001101010100",
		b"000000000111001001100111",
		b"000000000111000101101010",
		b"000000000111000001011111",
		b"000000000110111101000100",
		b"000000000110111000011100",
		b"000000000110110011100101",
		b"000000000110101110100001",
		b"000000000110101001001110",
		b"000000000110100011101110",
		b"000000000110011110000001",
		b"000000000110011000000110",
		b"000000000110010001111111",
		b"000000000110001011101011",
		b"000000000110000101001011",
		b"000000000101111110011111",
		b"000000000101110111101000",
		b"000000000101110000100100",
		b"000000000101101001010110",
		b"000000000101100001111100",
		b"000000000101011010011000",
		b"000000000101010010101010",
		b"000000000101001010110010",
		b"000000000101000010101111",
		b"000000000100111010100100",
		b"000000000100110010001111",
		b"000000000100101001110010",
		b"000000000100100001001100",
		b"000000000100011000011111",
		b"000000000100001111101001",
		b"000000000100000110101100",
		b"000000000011111101101000",
		b"000000000011110100011101",
		b"000000000011101011001011",
		b"000000000011100001110100",
		b"000000000011011000010110",
		b"000000000011001110110100",
		b"000000000011000101001100",
		b"000000000010111011011111",
		b"000000000010110001101111",
		b"000000000010100111111010",
		b"000000000010011110000001",
		b"000000000010010100000101",
		b"000000000010001010000111",
		b"000000000010000000000101",
		b"000000000001110110000010",
		b"000000000001101011111100",
		b"000000000001100001110110",
		b"000000000001010111101101",
		b"000000000001001101100100",
		b"000000000001000011011011",
		b"000000000000111001010001",
		b"000000000000101111001000",
		b"000000000000100100111111",
		b"000000000000011010111000",
		b"000000000000010000110001",
		b"000000000000000110101100",
		b"111111111111111100101001",
		b"111111111111110010101001",
		b"111111111111101000101011",
		b"111111111111011110110000",
		b"111111111111010100111000",
		b"111111111111001011000100",
		b"111111111111000001010100",
		b"111111111110110111101000",
		b"111111111110101110000001",
		b"111111111110100100011110",
		b"111111111110011011000001",
		b"111111111110010001101010",
		b"111111111110001000011000",
		b"111111111101111111001100",
		b"111111111101110110000111",
		b"111111111101101101001000",
		b"111111111101100100010001",
		b"111111111101011011100001",
		b"111111111101010010111000",
		b"111111111101001010010111",
		b"111111111101000001111111",
		b"111111111100111001101110",
		b"111111111100110001100111",
		b"111111111100101001101000",
		b"111111111100100001110010",
		b"111111111100011010000101",
		b"111111111100010010100011",
		b"111111111100001011001001",
		b"111111111100000011111010",
		b"111111111011111100110110",
		b"111111111011110101111011",
		b"111111111011101111001011",
		b"111111111011101000100111",
		b"111111111011100010001101",
		b"111111111011011011111110",
		b"111111111011010101111011",
		b"111111111011010000000011",
		b"111111111011001010010111",
		b"111111111011000100110111",
		b"111111111010111111100010",
		b"111111111010111010011010",
		b"111111111010110101011111",
		b"111111111010110000101111",
		b"111111111010101100001101",
		b"111111111010100111110110",
		b"111111111010100011101101",
		b"111111111010011111110000",
		b"111111111010011100000001",
		b"111111111010011000011110",
		b"111111111010010101001000",
		b"111111111010010010000000",
		b"111111111010001111000101",
		b"111111111010001100010111",
		b"111111111010001001110110",
		b"111111111010000111100011",
		b"111111111010000101011101",
		b"111111111010000011100101",
		b"111111111010000001111010",
		b"111111111010000000011100",
		b"111111111001111111001100",
		b"111111111001111110001001",
		b"111111111001111101010100",
		b"111111111001111100101100",
		b"111111111001111100010001",
		b"111111111001111100000100",
		b"111111111001111100000100",
		b"111111111001111100010010",
		b"111111111001111100101100",
		b"111111111001111101010100",
		b"111111111001111110001001",
		b"111111111001111111001011",
		b"111111111010000000011001",
		b"111111111010000001110101",
		b"111111111010000011011101",
		b"111111111010000101010010",
		b"111111111010000111010100",
		b"111111111010001001100001",
		b"111111111010001011111100",
		b"111111111010001110100010",
		b"111111111010010001010100",
		b"111111111010010100010010",
		b"111111111010010111011100",
		b"111111111010011010110010",
		b"111111111010011110010011",
		b"111111111010100001111111",
		b"111111111010100101110110",
		b"111111111010101001111001",
		b"111111111010101110000110",
		b"111111111010110010011101",
		b"111111111010110110111111",
		b"111111111010111011101100",
		b"111111111011000000100010",
		b"111111111011000101100010",
		b"111111111011001010101011",
		b"111111111011001111111110",
		b"111111111011010101011010",
		b"111111111011011010111111",
		b"111111111011100000101101",
		b"111111111011100110100100",
		b"111111111011101100100010",
		b"111111111011110010101001",
		b"111111111011111000110111",
		b"111111111011111111001101",
		b"111111111100000101101010",
		b"111111111100001100001110",
		b"111111111100010010111001",
		b"111111111100011001101011",
		b"111111111100100000100011",
		b"111111111100100111100001",
		b"111111111100101110100100",
		b"111111111100110101101110",
		b"111111111100111100111100",
		b"111111111101000100001111",
		b"111111111101001011101000",
		b"111111111101010011000100",
		b"111111111101011010100101",
		b"111111111101100010001010",
		b"111111111101101001110010",
		b"111111111101110001011110",
		b"111111111101111001001100",
		b"111111111110000000111110",
		b"111111111110001000110010",
		b"111111111110010000101000",
		b"111111111110011000100000",
		b"111111111110100000011010",
		b"111111111110101000010101",
		b"111111111110110000010010",
		b"111111111110111000001111",
		b"111111111111000000001101",
		b"111111111111001000001011",
		b"111111111111010000001010",
		b"111111111111011000001000",
		b"111111111111100000000101",
		b"111111111111101000000010",
		b"111111111111101111111110",
		b"111111111111110111111000",
		b"111111111111111111110001",
		b"000000000000000111101000",
		b"000000000000001111011100",
		b"000000000000010111001111",
		b"000000000000011110111111",
		b"000000000000100110101011",
		b"000000000000101110010101",
		b"000000000000110101111100",
		b"000000000000111101011110",
		b"000000000001000100111101",
		b"000000000001001100011000",
		b"000000000001010011101110",
		b"000000000001011011000000",
		b"000000000001100010001101",
		b"000000000001101001010101",
		b"000000000001110000011000",
		b"000000000001110111010101",
		b"000000000001111110001100",
		b"000000000010000100111101",
		b"000000000010001011101001",
		b"000000000010010010001110",
		b"000000000010011000101100",
		b"000000000010011111000011",
		b"000000000010100101010100",
		b"000000000010101011011110",
		b"000000000010110001100000",
		b"000000000010110111011010",
		b"000000000010111101001101",
		b"000000000011000010111001",
		b"000000000011001000011100",
		b"000000000011001101110111",
		b"000000000011010011001001",
		b"000000000011011000010011",
		b"000000000011011101010101",
		b"000000000011100010001101",
		b"000000000011100110111101",
		b"000000000011101011100100",
		b"000000000011110000000010",
		b"000000000011110100010110",
		b"000000000011111000100001",
		b"000000000011111100100010",
		b"000000000100000000011010",
		b"000000000100000100001000",
		b"000000000100000111101101",
		b"000000000100001011000111",
		b"000000000100001110010111",
		b"000000000100010001011110",
		b"000000000100010100011010",
		b"000000000100010111001100",
		b"000000000100011001110100",
		b"000000000100011100010010",
		b"000000000100011110100101",
		b"000000000100100000101110",
		b"000000000100100010101101",
		b"000000000100100100100001",
		b"000000000100100110001010",
		b"000000000100100111101001",
		b"000000000100101000111110",
		b"000000000100101010001000",
		b"000000000100101011001000",
		b"000000000100101011111101",
		b"000000000100101100100111",
		b"000000000100101101000111",
		b"000000000100101101011101",
		b"000000000100101101101000",
		b"000000000100101101101001",
		b"000000000100101101100000",
		b"000000000100101101001100",
		b"000000000100101100101110",
		b"000000000100101100000101",
		b"000000000100101011010011",
		b"000000000100101010010110",
		b"000000000100101001010000",
		b"000000000100100111111111",
		b"000000000100100110100101",
		b"000000000100100101000000",
		b"000000000100100011010010",
		b"000000000100100001011011",
		b"000000000100011111011010",
		b"000000000100011101001111",
		b"000000000100011010111011",
		b"000000000100011000011110",
		b"000000000100010101111000",
		b"000000000100010011001001",
		b"000000000100010000010001",
		b"000000000100001101010001",
		b"000000000100001010001000",
		b"000000000100000110110110",
		b"000000000100000011011100",
		b"000000000011111111111010",
		b"000000000011111100010000",
		b"000000000011111000011110",
		b"000000000011110100100101",
		b"000000000011110000100100",
		b"000000000011101100011011",
		b"000000000011101000001011",
		b"000000000011100011110101",
		b"000000000011011111010111",
		b"000000000011011010110011",
		b"000000000011010110001000",
		b"000000000011010001010111",
		b"000000000011001100100000",
		b"000000000011000111100011",
		b"000000000011000010100000",
		b"000000000010111101011000",
		b"000000000010111000001010",
		b"000000000010110010110111",
		b"000000000010101101011111",
		b"000000000010101000000010",
		b"000000000010100010100001",
		b"000000000010011100111011",
		b"000000000010010111010001",
		b"000000000010010001100100",
		b"000000000010001011110010",
		b"000000000010000101111101",
		b"000000000010000000000100",
		b"000000000001111010001001",
		b"000000000001110100001010",
		b"000000000001101110001001",
		b"000000000001101000000101",
		b"000000000001100001111111",
		b"000000000001011011110111",
		b"000000000001010101101110",
		b"000000000001001111100010",
		b"000000000001001001010101",
		b"000000000001000011000111",
		b"000000000000111100111000",
		b"000000000000110110101000",
		b"000000000000110000011000",
		b"000000000000101010000111",
		b"000000000000100011110110",
		b"000000000000011101100101",
		b"000000000000010111010101",
		b"000000000000010001000101",
		b"000000000000001010110101",
		b"000000000000000100100111",
		b"111111111111111110011001",
		b"111111111111111000001110",
		b"111111111111110010000011",
		b"111111111111101011111010",
		b"111111111111100101110100",
		b"111111111111011111101111",
		b"111111111111011001101101",
		b"111111111111010011101101",
		b"111111111111001101110000",
		b"111111111111000111110110",
		b"111111111111000001111111",
		b"111111111110111100001011",
		b"111111111110110110011011",
		b"111111111110110000101110",
		b"111111111110101011000110",
		b"111111111110100101100001",
		b"111111111110100000000000",
		b"111111111110011010100100",
		b"111111111110010101001100",
		b"111111111110001111111001",
		b"111111111110001010101011",
		b"111111111110000101100010",
		b"111111111110000000011110",
		b"111111111101111011011111",
		b"111111111101110110100110",
		b"111111111101110001110010",
		b"111111111101101101000100",
		b"111111111101101000011100",
		b"111111111101100011111010",
		b"111111111101011111011110",
		b"111111111101011011001000",
		b"111111111101010110111001",
		b"111111111101010010110000",
		b"111111111101001110101110",
		b"111111111101001010110011",
		b"111111111101000110111110",
		b"111111111101000011010001",
		b"111111111100111111101010",
		b"111111111100111100001011",
		b"111111111100111000110011",
		b"111111111100110101100010",
		b"111111111100110010011000",
		b"111111111100101111010110",
		b"111111111100101100011100",
		b"111111111100101001101001",
		b"111111111100100110111110",
		b"111111111100100100011011",
		b"111111111100100001111111",
		b"111111111100011111101100",
		b"111111111100011101100000",
		b"111111111100011011011100",
		b"111111111100011001100000",
		b"111111111100010111101101",
		b"111111111100010110000001",
		b"111111111100010100011101",
		b"111111111100010011000010",
		b"111111111100010001101110",
		b"111111111100010000100011",
		b"111111111100001111100000",
		b"111111111100001110100101",
		b"111111111100001101110010",
		b"111111111100001101001000",
		b"111111111100001100100101",
		b"111111111100001100001011",
		b"111111111100001011111000",
		b"111111111100001011101110",
		b"111111111100001011101100",
		b"111111111100001011110010",
		b"111111111100001100000000",
		b"111111111100001100010110",
		b"111111111100001100110100",
		b"111111111100001101011001",
		b"111111111100001110000111",
		b"111111111100001110111100",
		b"111111111100001111111001",
		b"111111111100010000111110",
		b"111111111100010010001010",
		b"111111111100010011011110",
		b"111111111100010100111001",
		b"111111111100010110011100",
		b"111111111100011000000110",
		b"111111111100011001110111",
		b"111111111100011011110000",
		b"111111111100011101101111",
		b"111111111100011111110101",
		b"111111111100100010000010",
		b"111111111100100100010110",
		b"111111111100100110110001",
		b"111111111100101001010010",
		b"111111111100101011111001",
		b"111111111100101110100111",
		b"111111111100110001011011",
		b"111111111100110100010101",
		b"111111111100110111010101",
		b"111111111100111010011011",
		b"111111111100111101100111",
		b"111111111101000000111000",
		b"111111111101000100001111",
		b"111111111101000111101011",
		b"111111111101001011001100",
		b"111111111101001110110010",
		b"111111111101010010011110",
		b"111111111101010110001110",
		b"111111111101011010000010",
		b"111111111101011101111011",
		b"111111111101100001111000",
		b"111111111101100101111010",
		b"111111111101101010000000",
		b"111111111101101110001001",
		b"111111111101110010010110",
		b"111111111101110110100111",
		b"111111111101111010111011",
		b"111111111101111111010011",
		b"111111111110000011101101",
		b"111111111110001000001011",
		b"111111111110001100101011",
		b"111111111110010001001110",
		b"111111111110010101110011",
		b"111111111110011010011010",
		b"111111111110011111000100",
		b"111111111110100011110000",
		b"111111111110101000011101",
		b"111111111110101101001100",
		b"111111111110110001111101",
		b"111111111110110110101111",
		b"111111111110111011100010",
		b"111111111111000000010101",
		b"111111111111000101001010",
		b"111111111111001010000000",
		b"111111111111001110110101",
		b"111111111111010011101100",
		b"111111111111011000100010",
		b"111111111111011101011000",
		b"111111111111100010001110",
		b"111111111111100111000100",
		b"111111111111101011111001",
		b"111111111111110000101110",
		b"111111111111110101100001",
		b"111111111111111010010100",
		b"111111111111111111000101",
		b"000000000000000011110110",
		b"000000000000001000100101",
		b"000000000000001101010010",
		b"000000000000010001111101",
		b"000000000000010110100111",
		b"000000000000011011001110",
		b"000000000000011111110011",
		b"000000000000100100010110",
		b"000000000000101000110111",
		b"000000000000101101010100",
		b"000000000000110001101111",
		b"000000000000110110000111",
		b"000000000000111010011100",
		b"000000000000111110101110",
		b"000000000001000010111100",
		b"000000000001000111000111",
		b"000000000001001011001110",
		b"000000000001001111010010",
		b"000000000001010011010010",
		b"000000000001010111001110",
		b"000000000001011011000101",
		b"000000000001011110111001",
		b"000000000001100010101000",
		b"000000000001100110010011",
		b"000000000001101001111001",
		b"000000000001101101011011",
		b"000000000001110000111000",
		b"000000000001110100010000",
		b"000000000001110111100011",
		b"000000000001111010110001",
		b"000000000001111101111010",
		b"000000000010000000111110",
		b"000000000010000011111101",
		b"000000000010000110110110",
		b"000000000010001001101010",
		b"000000000010001100011000",
		b"000000000010001111000000",
		b"000000000010010001100011",
		b"000000000010010100000000",
		b"000000000010010110011000",
		b"000000000010011000101001",
		b"000000000010011010110101",
		b"000000000010011100111011",
		b"000000000010011110111010",
		b"000000000010100000110100",
		b"000000000010100010100111",
		b"000000000010100100010101",
		b"000000000010100101111100",
		b"000000000010100111011101",
		b"000000000010101000110111",
		b"000000000010101010001100",
		b"000000000010101011011010",
		b"000000000010101100100010",
		b"000000000010101101100011",
		b"000000000010101110011110",
		b"000000000010101111010011",
		b"000000000010110000000001",
		b"000000000010110000101001",
		b"000000000010110001001011",
		b"000000000010110001100110",
		b"000000000010110001111011",
		b"000000000010110010001001",
		b"000000000010110010010001",
		b"000000000010110010010011",
		b"000000000010110010001111",
		b"000000000010110010000100",
		b"000000000010110001110011",
		b"000000000010110001011100",
		b"000000000010110000111110",
		b"000000000010110000011011",
		b"000000000010101111110001",
		b"000000000010101111000001",
		b"000000000010101110001011",
		b"000000000010101101001111",
		b"000000000010101100001110",
		b"000000000010101011000110",
		b"000000000010101001111000",
		b"000000000010101000100101",
		b"000000000010100111001100",
		b"000000000010100101101101",
		b"000000000010100100001001",
		b"000000000010100010011111",
		b"000000000010100000110000",
		b"000000000010011110111011",
		b"000000000010011101000001",
		b"000000000010011011000010",
		b"000000000010011000111101",
		b"000000000010010110110100",
		b"000000000010010100100101",
		b"000000000010010010010010",
		b"000000000010001111111010",
		b"000000000010001101011101",
		b"000000000010001010111100",
		b"000000000010001000010110",
		b"000000000010000101101011",
		b"000000000010000010111101",
		b"000000000010000000001010",
		b"000000000001111101010011",
		b"000000000001111010011000",
		b"000000000001110111011001",
		b"000000000001110100010110",
		b"000000000001110001001111",
		b"000000000001101110000101",
		b"000000000001101010111000",
		b"000000000001100111100111",
		b"000000000001100100010011",
		b"000000000001100000111100",
		b"000000000001011101100010",
		b"000000000001011010000101",
		b"000000000001010110100101",
		b"000000000001010011000011",
		b"000000000001001111011110",
		b"000000000001001011110110",
		b"000000000001001000001101",
		b"000000000001000100100001",
		b"000000000001000000110011",
		b"000000000000111101000100",
		b"000000000000111001010010",
		b"000000000000110101011111",
		b"000000000000110001101011",
		b"000000000000101101110101",
		b"000000000000101001111101",
		b"000000000000100110000101",
		b"000000000000100010001100",
		b"000000000000011110010001",
		b"000000000000011010010110",
		b"000000000000010110011011",
		b"000000000000010010011111",
		b"000000000000001110100010",
		b"000000000000001010100110",
		b"000000000000000110101001",
		b"000000000000000010101100",
		b"111111111111111110101111",
		b"111111111111111010110011",
		b"111111111111110110110111",
		b"111111111111110010111011",
		b"111111111111101111000001",
		b"111111111111101011000110",
		b"111111111111100111001101",
		b"111111111111100011010101",
		b"111111111111011111011110",
		b"111111111111011011101000",
		b"111111111111010111110100",
		b"111111111111010100000001",
		b"111111111111010000001111",
		b"111111111111001100011111",
		b"111111111111001000110001",
		b"111111111111000101000110",
		b"111111111111000001011100",
		b"111111111110111101110100",
		b"111111111110111010001110",
		b"111111111110110110101011",
		b"111111111110110011001010",
		b"111111111110101111101100",
		b"111111111110101100010001",
		b"111111111110101000111000",
		b"111111111110100101100010",
		b"111111111110100010001111",
		b"111111111110011111000000",
		b"111111111110011011110011",
		b"111111111110011000101001",
		b"111111111110010101100011",
		b"111111111110010010100001",
		b"111111111110001111100001",
		b"111111111110001100100110",
		b"111111111110001001101110",
		b"111111111110000110111010",
		b"111111111110000100001001",
		b"111111111110000001011101",
		b"111111111101111110110100",
		b"111111111101111100010000",
		b"111111111101111001101111",
		b"111111111101110111010011",
		b"111111111101110100111011",
		b"111111111101110010101000",
		b"111111111101110000011000",
		b"111111111101101110001101",
		b"111111111101101100000111",
		b"111111111101101010000101",
		b"111111111101101000000111",
		b"111111111101100110001110",
		b"111111111101100100011010",
		b"111111111101100010101010",
		b"111111111101100001000000",
		b"111111111101011111011001",
		b"111111111101011101111000",
		b"111111111101011100011100",
		b"111111111101011011000100",
		b"111111111101011001110001",
		b"111111111101011000100011",
		b"111111111101010111011010",
		b"111111111101010110010110",
		b"111111111101010101010111",
		b"111111111101010100011101",
		b"111111111101010011101000",
		b"111111111101010010111000",
		b"111111111101010010001101",
		b"111111111101010001100111",
		b"111111111101010001000101",
		b"111111111101010000101001",
		b"111111111101010000010010",
		b"111111111101010000000000",
		b"111111111101001111110011",
		b"111111111101001111101010",
		b"111111111101001111100111",
		b"111111111101001111101001",
		b"111111111101001111101111",
		b"111111111101001111111011",
		b"111111111101010000001011",
		b"111111111101010000100000",
		b"111111111101010000111010",
		b"111111111101010001011001",
		b"111111111101010001111100",
		b"111111111101010010100100",
		b"111111111101010011010001",
		b"111111111101010100000010",
		b"111111111101010100111000",
		b"111111111101010101110011",
		b"111111111101010110110010",
		b"111111111101010111110110",
		b"111111111101011000111110",
		b"111111111101011010001010",
		b"111111111101011011011011",
		b"111111111101011100110000",
		b"111111111101011110001001",
		b"111111111101011111100110",
		b"111111111101100001000111",
		b"111111111101100010101101",
		b"111111111101100100010110",
		b"111111111101100110000011",
		b"111111111101100111110100",
		b"111111111101101001101000",
		b"111111111101101011100001",
		b"111111111101101101011101",
		b"111111111101101111011100",
		b"111111111101110001011111",
		b"111111111101110011100101",
		b"111111111101110101101111",
		b"111111111101110111111011",
		b"111111111101111010001011",
		b"111111111101111100011110",
		b"111111111101111110110100",
		b"111111111110000001001101",
		b"111111111110000011101000",
		b"111111111110000110000110",
		b"111111111110001000100111",
		b"111111111110001011001010",
		b"111111111110001101110000",
		b"111111111110010000011000",
		b"111111111110010011000010",
		b"111111111110010101101111",
		b"111111111110011000011101",
		b"111111111110011011001101",
		b"111111111110011110000000",
		b"111111111110100000110100",
		b"111111111110100011101001",
		b"111111111110100110100001",
		b"111111111110101001011010",
		b"111111111110101100010100",
		b"111111111110101111001111",
		b"111111111110110010001100",
		b"111111111110110101001001",
		b"111111111110111000001000",
		b"111111111110111011001000",
		b"111111111110111110001000",
		b"111111111111000001001001",
		b"111111111111000100001011",
		b"111111111111000111001101",
		b"111111111111001010001111",
		b"111111111111001101010010",
		b"111111111111010000010101",
		b"111111111111010011011000",
		b"111111111111010110011011",
		b"111111111111011001011110",
		b"111111111111011100100000",
		b"111111111111011111100011",
		b"111111111111100010100101",
		b"111111111111100101100110",
		b"111111111111101000100111",
		b"111111111111101011100111",
		b"111111111111101110100111",
		b"111111111111110001100101",
		b"111111111111110100100011",
		b"111111111111110111011111",
		b"111111111111111010011010",
		b"111111111111111101010100",
		b"000000000000000000001101",
		b"000000000000000011000100",
		b"000000000000000101111010",
		b"000000000000001000101110",
		b"000000000000001011100000",
		b"000000000000001110010001",
		b"000000000000010001000000",
		b"000000000000010011101100",
		b"000000000000010110010111",
		b"000000000000011001000000",
		b"000000000000011011100110",
		b"000000000000011110001010",
		b"000000000000100000101100",
		b"000000000000100011001011",
		b"000000000000100101101000",
		b"000000000000101000000010",
		b"000000000000101010011001",
		b"000000000000101100101110",
		b"000000000000101111000000",
		b"000000000000110001001111",
		b"000000000000110011011011",
		b"000000000000110101100101",
		b"000000000000110111101011",
		b"000000000000111001101110",
		b"000000000000111011101101",
		b"000000000000111101101010",
		b"000000000000111111100011",
		b"000000000001000001011001",
		b"000000000001000011001011",
		b"000000000001000100111010",
		b"000000000001000110100110",
		b"000000000001001000001110",
		b"000000000001001001110010",
		b"000000000001001011010010",
		b"000000000001001100101111",
		b"000000000001001110001000",
		b"000000000001001111011110",
		b"000000000001010000101111",
		b"000000000001010001111101",
		b"000000000001010011000111",
		b"000000000001010100001101",
		b"000000000001010101001110",
		b"000000000001010110001100",
		b"000000000001010111000110",
		b"000000000001010111111100",
		b"000000000001011000101110",
		b"000000000001011001011011",
		b"000000000001011010000101",
		b"000000000001011010101010",
		b"000000000001011011001011",
		b"000000000001011011101000",
		b"000000000001011100000001",
		b"000000000001011100010110",
		b"000000000001011100100111",
		b"000000000001011100110011",
		b"000000000001011100111011",
		b"000000000001011100111111",
		b"000000000001011100111111",
		b"000000000001011100111010",
		b"000000000001011100110010",
		b"000000000001011100100101",
		b"000000000001011100010100",
		b"000000000001011011111111",
		b"000000000001011011100101",
		b"000000000001011011001000",
		b"000000000001011010100110",
		b"000000000001011010000000",
		b"000000000001011001010110",
		b"000000000001011000101000",
		b"000000000001010111110110",
		b"000000000001010111000000",
		b"000000000001010110000101",
		b"000000000001010101000111",
		b"000000000001010100000101",
		b"000000000001010010111111",
		b"000000000001010001110100",
		b"000000000001010000100110",
		b"000000000001001111010101",
		b"000000000001001101111111",
		b"000000000001001100100101",
		b"000000000001001011001000",
		b"000000000001001001100111",
		b"000000000001001000000011",
		b"000000000001000110011010",
		b"000000000001000100101111",
		b"000000000001000010111111",
		b"000000000001000001001100",
		b"000000000000111111010110",
		b"000000000000111101011100",
		b"000000000000111011011111",
		b"000000000000111001011111",
		b"000000000000110111011011",
		b"000000000000110101010101",
		b"000000000000110011001011",
		b"000000000000110000111110",
		b"000000000000101110101110",
		b"000000000000101100011011",
		b"000000000000101010000101",
		b"000000000000100111101101",
		b"000000000000100101010001",
		b"000000000000100010110011",
		b"000000000000100000010010",
		b"000000000000011101101111",
		b"000000000000011011001001",
		b"000000000000011000100000",
		b"000000000000010101110110",
		b"000000000000010011001001",
		b"000000000000010000011001",
		b"000000000000001101101000",
		b"000000000000001010110100",
		b"000000000000000111111111",
		b"000000000000000101000111",
		b"000000000000000010001101",
		b"111111111111111111010010",
		b"111111111111111100010101",
		b"111111111111111001010110",
		b"111111111111110110010110",
		b"111111111111110011010100",
		b"111111111111110000010000",
		b"111111111111101101001100",
		b"111111111111101010000110",
		b"111111111111100110111110",
		b"111111111111100011110110",
		b"111111111111100000101100",
		b"111111111111011101100010",
		b"111111111111011010010110",
		b"111111111111010111001010",
		b"111111111111010011111101",
		b"111111111111010000101111",
		b"111111111111001101100001",
		b"111111111111001010010010",
		b"111111111111000111000010",
		b"111111111111000011110010",
		b"111111111111000000100010",
		b"111111111110111101010010",
		b"111111111110111010000001",
		b"111111111110110110110001",
		b"111111111110110011100000",
		b"111111111110110000010000",
		b"111111111110101100111111",
		b"111111111110101001101111",
		b"111111111110100110011111",
		b"111111111110100011001111",
		b"111111111110100000000000",
		b"111111111110011100110010",
		b"111111111110011001100100",
		b"111111111110010110010110",
		b"111111111110010011001001",
		b"111111111110001111111110",
		b"111111111110001100110011",
		b"111111111110001001101001",
		b"111111111110000110011111",
		b"111111111110000011010111",
		b"111111111110000000010001",
		b"111111111101111101001011",
		b"111111111101111010000111",
		b"111111111101110111000100",
		b"111111111101110100000010",
		b"111111111101110001000010",
		b"111111111101101110000011",
		b"111111111101101011000110",
		b"111111111101101000001011",
		b"111111111101100101010010",
		b"111111111101100010011010",
		b"111111111101011111100100",
		b"111111111101011100110000",
		b"111111111101011001111110",
		b"111111111101010111001110",
		b"111111111101010100100000",
		b"111111111101010001110100",
		b"111111111101001111001010",
		b"111111111101001100100011",
		b"111111111101001001111110",
		b"111111111101000111011011",
		b"111111111101000100111010",
		b"111111111101000010011100",
		b"111111111101000000000001",
		b"111111111100111101101000",
		b"111111111100111011010001",
		b"111111111100111000111110",
		b"111111111100110110101101",
		b"111111111100110100011110",
		b"111111111100110010010010",
		b"111111111100110000001010",
		b"111111111100101110000011",
		b"111111111100101100000000",
		b"111111111100101010000000",
		b"111111111100101000000011",
		b"111111111100100110001000",
		b"111111111100100100010001",
		b"111111111100100010011100",
		b"111111111100100000101011",
		b"111111111100011110111101",
		b"111111111100011101010001",
		b"111111111100011011101001",
		b"111111111100011010000101",
		b"111111111100011000100011",
		b"111111111100010111000100",
		b"111111111100010101101001",
		b"111111111100010100010001",
		b"111111111100010010111100",
		b"111111111100010001101011",
		b"111111111100010000011101",
		b"111111111100001111010010",
		b"111111111100001110001010",
		b"111111111100001101000110",
		b"111111111100001100000101",
		b"111111111100001011001000",
		b"111111111100001010001110",
		b"111111111100001001010111",
		b"111111111100001000100100",
		b"111111111100000111110100",
		b"111111111100000111000111",
		b"111111111100000110011110",
		b"111111111100000101111000",
		b"111111111100000101010110",
		b"111111111100000100110111",
		b"111111111100000100011011",
		b"111111111100000100000011",
		b"111111111100000011101110",
		b"111111111100000011011100",
		b"111111111100000011001110",
		b"111111111100000011000100",
		b"111111111100000010111100",
		b"111111111100000010111000",
		b"111111111100000010110111",
		b"111111111100000010111010",
		b"111111111100000011000000",
		b"111111111100000011001001",
		b"111111111100000011010110",
		b"111111111100000011100101",
		b"111111111100000011111000",
		b"111111111100000100001110",
		b"111111111100000100101000",
		b"111111111100000101000100",
		b"111111111100000101100100",
		b"111111111100000110000111",
		b"111111111100000110101101",
		b"111111111100000111010110",
		b"111111111100001000000010",
		b"111111111100001000110010",
		b"111111111100001001100100",
		b"111111111100001010011001",
		b"111111111100001011010001",
		b"111111111100001100001100",
		b"111111111100001101001010",
		b"111111111100001110001011",
		b"111111111100001111001111",
		b"111111111100010000010101",
		b"111111111100010001011110",
		b"111111111100010010101010",
		b"111111111100010011111001",
		b"111111111100010101001010",
		b"111111111100010110011110",
		b"111111111100010111110101",
		b"111111111100011001001110",
		b"111111111100011010101010",
		b"111111111100011100001000",
		b"111111111100011101101000",
		b"111111111100011111001011",
		b"111111111100100000110000",
		b"111111111100100010011000",
		b"111111111100100100000010",
		b"111111111100100101101110",
		b"111111111100100111011100",
		b"111111111100101001001101",
		b"111111111100101010111111",
		b"111111111100101100110100",
		b"111111111100101110101010",
		b"111111111100110000100011",
		b"111111111100110010011110",
		b"111111111100110100011010",
		b"111111111100110110011000",
		b"111111111100111000011000",
		b"111111111100111010011010",
		b"111111111100111100011110",
		b"111111111100111110100011",
		b"111111111101000000101010",
		b"111111111101000010110010",
		b"111111111101000100111100",
		b"111111111101000111000111",
		b"111111111101001001010100",
		b"111111111101001011100010",
		b"111111111101001101110001",
		b"111111111101010000000010",
		b"111111111101010010010100",
		b"111111111101010100100111",
		b"111111111101010110111100",
		b"111111111101011001010001",
		b"111111111101011011100111",
		b"111111111101011101111111",
		b"111111111101100000010111",
		b"111111111101100010110000",
		b"111111111101100101001011",
		b"111111111101100111100110",
		b"111111111101101010000001",
		b"111111111101101100011110",
		b"111111111101101110111011",
		b"111111111101110001011001",
		b"111111111101110011110111",
		b"111111111101110110010110",
		b"111111111101111000110101",
		b"111111111101111011010101",
		b"111111111101111101110101",
		b"111111111110000000010101",
		b"111111111110000010110110",
		b"111111111110000101010111",
		b"111111111110000111111001",
		b"111111111110001010011010",
		b"111111111110001100111100",
		b"111111111110001111011101",
		b"111111111110010001111111",
		b"111111111110010100100001",
		b"111111111110010111000010",
		b"111111111110011001100100",
		b"111111111110011100000101",
		b"111111111110011110100110",
		b"111111111110100001001000",
		b"111111111110100011101000",
		b"111111111110100110001001",
		b"111111111110101000101001",
		b"111111111110101011001001",
		b"111111111110101101101000",
		b"111111111110110000000111",
		b"111111111110110010100110",
		b"111111111110110101000100",
		b"111111111110110111100001",
		b"111111111110111001111110",
		b"111111111110111100011010",
		b"111111111110111110110101",
		b"111111111111000001010000",
		b"111111111111000011101010",
		b"111111111111000110000100",
		b"111111111111001000011100",
		b"111111111111001010110100",
		b"111111111111001101001011",
		b"111111111111001111100001",
		b"111111111111010001110110",
		b"111111111111010100001010",
		b"111111111111010110011101",
		b"111111111111011000101111",
		b"111111111111011011000000",
		b"111111111111011101010000",
		b"111111111111011111011111",
		b"111111111111100001101101",
		b"111111111111100011111001",
		b"111111111111100110000101",
		b"111111111111101000001111",
		b"111111111111101010011000",
		b"111111111111101100100000",
		b"111111111111101110100110",
		b"111111111111110000101011",
		b"111111111111110010101111",
		b"111111111111110100110010",
		b"111111111111110110110011",
		b"111111111111111000110011",
		b"111111111111111010110010",
		b"111111111111111100101111",
		b"111111111111111110101010",
		b"000000000000000000100100",
		b"000000000000000010011101",
		b"000000000000000100010101",
		b"000000000000000110001010",
		b"000000000000000111111111",
		b"000000000000001001110001",
		b"000000000000001011100011",
		b"000000000000001101010010",
		b"000000000000001111000001",
		b"000000000000010000101101",
		b"000000000000010010011000",
		b"000000000000010100000010",
		b"000000000000010101101010",
		b"000000000000010111010000",
		b"000000000000011000110101",
		b"000000000000011010011000",
		b"000000000000011011111001",
		b"000000000000011101011001",
		b"000000000000011110110111",
		b"000000000000100000010011",
		b"000000000000100001101110",
		b"000000000000100011000111",
		b"000000000000100100011111",
		b"000000000000100101110101",
		b"000000000000100111001001",
		b"000000000000101000011100",
		b"000000000000101001101101",
		b"000000000000101010111100",
		b"000000000000101100001001",
		b"000000000000101101010101",
		b"000000000000101110100000",
		b"000000000000101111101000",
		b"000000000000110000101111",
		b"000000000000110001110100",
		b"000000000000110010111000",
		b"000000000000110011111010",
		b"000000000000110100111010",
		b"000000000000110101111001",
		b"000000000000110110110110",
		b"000000000000110111110001",
		b"000000000000111000101011",
		b"000000000000111001100011",
		b"000000000000111010011010",
		b"000000000000111011001111",
		b"000000000000111100000010",
		b"000000000000111100110100",
		b"000000000000111101100100",
		b"000000000000111110010010",
		b"000000000000111110111111",
		b"000000000000111111101011",
		b"000000000001000000010101",
		b"000000000001000000111101",
		b"000000000001000001100100",
		b"000000000001000010001001",
		b"000000000001000010101101",
		b"000000000001000011001111",
		b"000000000001000011110000",
		b"000000000001000100001111",
		b"000000000001000100101101",
		b"000000000001000101001001",
		b"000000000001000101100100",
		b"000000000001000101111110",
		b"000000000001000110010110",
		b"000000000001000110101101",
		b"000000000001000111000010",
		b"000000000001000111010110",
		b"000000000001000111101001",
		b"000000000001000111111010",
		b"000000000001001000001010",
		b"000000000001001000011001",
		b"000000000001001000100110",
		b"000000000001001000110010",
		b"000000000001001000111101",
		b"000000000001001001000110",
		b"000000000001001001001111",
		b"000000000001001001010110",
		b"000000000001001001011100",
		b"000000000001001001100001",
		b"000000000001001001100100",
		b"000000000001001001100111",
		b"000000000001001001101000",
		b"000000000001001001101000",
		b"000000000001001001100111",
		b"000000000001001001100101",
		b"000000000001001001100010",
		b"000000000001001001011110",
		b"000000000001001001011001",
		b"000000000001001001010011",
		b"000000000001001001001100",
		b"000000000001001001000100",
		b"000000000001001000111011",
		b"000000000001001000110001",
		b"000000000001001000100110",
		b"000000000001001000011010",
		b"000000000001001000001101",
		b"000000000001001000000000",
		b"000000000001000111110001",
		b"000000000001000111100010",
		b"000000000001000111010010",
		b"000000000001000111000001",
		b"000000000001000110110000",
		b"000000000001000110011101",
		b"000000000001000110001010",
		b"000000000001000101110110",
		b"000000000001000101100010",
		b"000000000001000101001101",
		b"000000000001000100110111",
		b"000000000001000100100000",
		b"000000000001000100001001",
		b"000000000001000011110001",
		b"000000000001000011011001",
		b"000000000001000011000000",
		b"000000000001000010100110",
		b"000000000001000010001100",
		b"000000000001000001110001",
		b"000000000001000001010110",
		b"000000000001000000111011",
		b"000000000001000000011110",
		b"000000000001000000000010",
		b"000000000000111111100101",
		b"000000000000111111000111",
		b"000000000000111110101001",
		b"000000000000111110001011",
		b"000000000000111101101100",
		b"000000000000111101001101",
		b"000000000000111100101110",
		b"000000000000111100001110",
		b"000000000000111011101110",
		b"000000000000111011001101",
		b"000000000000111010101101",
		b"000000000000111010001100",
		b"000000000000111001101011",
		b"000000000000111001001001",
		b"000000000000111000100111",
		b"000000000000111000000101",
		b"000000000000110111100011",
		b"000000000000110111000001",
		b"000000000000110110011110",
		b"000000000000110101111100",
		b"000000000000110101011001",
		b"000000000000110100110110",
		b"000000000000110100010011",
		b"000000000000110011110000",
		b"000000000000110011001100",
		b"000000000000110010101001",
		b"000000000000110010000101",
		b"000000000000110001100010",
		b"000000000000110000111110",
		b"000000000000110000011010",
		b"000000000000101111110111",
		b"000000000000101111010011",
		b"000000000000101110101111",
		b"000000000000101110001100",
		b"000000000000101101101000",
		b"000000000000101101000100",
		b"000000000000101100100001",
		b"000000000000101011111101",
		b"000000000000101011011010",
		b"000000000000101010110110",
		b"000000000000101010010011",
		b"000000000000101001101111",
		b"000000000000101001001100",
		b"000000000000101000101001",
		b"000000000000101000000110",
		b"000000000000100111100011",
		b"000000000000100111000000",
		b"000000000000100110011110",
		b"000000000000100101111011",
		b"000000000000100101011001",
		b"000000000000100100110111",
		b"000000000000100100010100",
		b"000000000000100011110011",
		b"000000000000100011010001",
		b"000000000000100010101111",
		b"000000000000100010001110",
		b"000000000000100001101101",
		b"000000000000100001001100",
		b"000000000000100000101011",
		b"000000000000100000001011",
		b"000000000000011111101010",
		b"000000000000011111001010",
		b"000000000000011110101011",
		b"000000000000011110001011",
		b"000000000000011101101100",
		b"000000000000011101001100",
		b"000000000000011100101110",
		b"000000000000011100001111",
		b"000000000000011011110001",
		b"000000000000011011010010",
		b"000000000000011010110101",
		b"000000000000011010010111",
		b"000000000000011001111010",
		b"000000000000011001011101",
		b"000000000000011001000000",
		b"000000000000011000100011",
		b"000000000000011000000111",
		b"000000000000010111101011",
		b"000000000000010111010000",
		b"000000000000010110110100",
		b"000000000000010110011001",
		b"000000000000010101111111",
		b"000000000000010101100100",
		b"000000000000010101001010",
		b"000000000000010100110000",
		b"000000000000010100010110",
		b"000000000000010011111101",
		b"000000000000010011100100",
		b"000000000000010011001011",
		b"000000000000010010110011",
		b"000000000000010010011011",
		b"000000000000010010000011",
		b"000000000000010001101100",
		b"000000000000010001010101",
		b"000000000000010000111110",
		b"000000000000010000100111",
		b"000000000000010000010001",
		b"000000000000001111111011",
		b"000000000000001111100101",
		b"000000000000001111010000",
		b"000000000000001110111011",
		b"000000000000001110100110",
		b"000000000000001110010010",
		b"000000000000001101111110",
		b"000000000000001101101010",
		b"000000000000001101010110",
		b"000000000000001101000011",
		b"000000000000001100110000",
		b"000000000000001100011101",
		b"000000000000001100001011",
		b"000000000000001011111001",
		b"000000000000001011100111",
		b"000000000000001011010110",
		b"000000000000001011000101",
		b"000000000000001010110100",
		b"000000000000001010100011",
		b"000000000000001010010011",
		b"000000000000001010000011",
		b"000000000000001001110011",
		b"000000000000001001100011",
		b"000000000000001001010100",
		b"000000000000001001000101",
		b"000000000000001000110111",
		b"000000000000001000101000",
		b"000000000000001000011010",
		b"000000000000001000001100",
		b"000000000000000111111111",
		b"000000000000000111110001",
		b"000000000000000111100100",
		b"000000000000000111010111",
		b"000000000000000111001011",
		b"000000000000000110111110",
		b"000000000000000110110010",
		b"000000000000000110100110",
		b"000000000000000110011011",
		b"000000000000000110001111",
		b"000000000000000110000100",
		b"000000000000000101111001",
		b"000000000000000101101111",
		b"000000000000000101100100",
		b"000000000000000101011010",
		b"000000000000000101010000",
		b"000000000000000101000110",
		b"000000000000000100111100",
		b"000000000000000100110011",
		b"000000000000000100101010",
		b"000000000000000100100001",
		b"000000000000000100011000",
		b"000000000000000100010000",
		b"000000000000000100000111",
		b"000000000000000011111111",
		b"000000000000000011110111",
		b"000000000000000011110000",
		b"000000000000000011101000",
		b"000000000000000011100001",
		b"000000000000000011011001",
		b"000000000000000011010010",
		b"000000000000000011001011",
		b"000000000000000011000101",
		b"000000000000000010111110",
		b"000000000000000010111000",
		b"000000000000000010110010",
		b"000000000000000010101100",
		b"000000000000000010100110",
		b"000000000000000010100000",
		b"000000000000000010011011",
		b"000000000000000010010101",
		b"000000000000000010010000",
		b"000000000000000010001011",
		b"000000000000000010000110",
		b"000000000000000010000001",
		b"000000000000000001111100",
		b"000000000000000001111000",
		b"000000000000000001110011",
		b"000000000000000001101111",
		b"000000000000000001101011",
		b"000000000000000001100111",
		b"000000000000000001100011",
		b"000000000000000001011111",
		b"000000000000000001011011",
		b"000000000000000001011000",
		b"000000000000000001010100",
		b"000000000000000001010001",
		b"000000000000000001001110",
		b"000000000000000001001010",
		b"000000000000000001000111",
		b"000000000000000001000100",
		b"000000000000000001000010",
		b"000000000000000000111111",
		b"000000000000000000111100",
		b"000000000000000000111010",
		b"000000000000000000110111",
		b"000000000000000000110101",
		b"000000000000000000110010",
		b"000000000000000000110000",
		b"000000000000000000101110",
		b"000000000000000000101100",
		b"000000000000000000101010",
		b"000000000000000000101000",
		b"000000000000000000100110",
		b"000000000000000000100100",
		b"000000000000000000100010",
		b"000000000000000000100001",
		b"000000000000000000011111",
		b"000000000000000000011110",
		b"000000000000000000011100",
		b"000000000000000000011011",
		b"000000000000000000011001",
		b"000000000000000000011000",
		b"000000000000000000010111",
		b"000000000000000000010101",
		b"000000000000000000010100",
		b"000000000000000000010011",
		b"000000000000000000010010",
		b"000000000000000000010001",
		b"000000000000000000010000",
		b"000000000000000000001111",
		b"000000000000000000001110",
		b"000000000000000000001101",
		b"000000000000000000001101",
		b"000000000000000000001100",
		b"000000000000000000001011",
		b"000000000000000000001010",
		b"000000000000000000001010",
		b"000000000000000000001001",
		b"000000000000000000001000",
		b"000000000000000000001000",
		b"000000000000000000000111",
		b"000000000000000000000111",
		b"000000000000000000000110",
		b"000000000000000000000110",
		b"000000000000000000000101",
		b"000000000000000000000101",
		b"000000000000000000000101",
		b"000000000000000000000100",
		b"000000000000000000000100",
		b"000000000000000000000100",
		b"000000000000000000000011",
		b"000000000000000000000011",
		b"000000000000000000000011",
		b"000000000000000000000010",
		b"000000000000000000000010",
		b"000000000000000000000010",
		b"000000000000000000000010",
		b"000000000000000000000010",
		b"000000000000000000000001",
		b"000000000000000000000001",
		b"000000000000000000000001",
		b"000000000000000000000001",
		b"000000000000000000000001",
		b"000000000000000000000001",
		b"000000000000000000000001",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000",
		b"000000000000000000000000"
	);

end src_rom_pkg;